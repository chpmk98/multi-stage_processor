
module adder_32 ( a, b, cin, sum, v );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output v;
  wire   n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318;

  AOI22_X4 U129 ( .A1(b[1]), .A2(a[1]), .B1(n161), .B2(n131), .ZN(n163) );
  OAI21_X4 U130 ( .B1(n159), .B2(n130), .A(n129), .ZN(n161) );
  OAI22_X4 U131 ( .A1(n136), .A2(n135), .B1(n167), .B2(n168), .ZN(n171) );
  NOR2_X2 U132 ( .A1(n187), .A2(n279), .ZN(n126) );
  AOI21_X2 U133 ( .B1(n101), .B2(n232), .A(n230), .ZN(n111) );
  NAND3_X2 U134 ( .A1(n256), .A2(n255), .A3(n118), .ZN(n264) );
  NOR2_X2 U135 ( .A1(n252), .A2(n212), .ZN(n117) );
  NAND3_X2 U136 ( .A1(n264), .A2(n263), .A3(n119), .ZN(n265) );
  NAND3_X2 U137 ( .A1(n207), .A2(n255), .A3(n256), .ZN(n119) );
  OAI21_X2 U138 ( .B1(n188), .B2(n97), .A(n282), .ZN(n190) );
  NOR3_X2 U139 ( .A1(n289), .A2(n291), .A3(n292), .ZN(n144) );
  NOR3_X2 U140 ( .A1(n300), .A2(n291), .A3(n292), .ZN(n107) );
  AOI21_X2 U141 ( .B1(n110), .B2(n238), .A(n109), .ZN(n112) );
  NOR2_X2 U142 ( .A1(n220), .A2(n230), .ZN(n110) );
  NOR2_X2 U143 ( .A1(n260), .A2(n201), .ZN(n120) );
  NAND3_X2 U144 ( .A1(n98), .A2(n271), .A3(n200), .ZN(n202) );
  NOR3_X2 U145 ( .A1(n152), .A2(n151), .A3(n150), .ZN(n153) );
  NAND3_X2 U146 ( .A1(n246), .A2(n245), .A3(n113), .ZN(n248) );
  NAND3_X2 U147 ( .A1(n254), .A2(n253), .A3(n116), .ZN(n255) );
  NAND3_X2 U148 ( .A1(n215), .A2(n248), .A3(n247), .ZN(n116) );
  OAI21_X2 U149 ( .B1(n189), .B2(n190), .A(n193), .ZN(n270) );
  NOR2_X2 U150 ( .A1(n185), .A2(n192), .ZN(n189) );
  NAND3_X2 U151 ( .A1(n205), .A2(n265), .A3(n266), .ZN(n122) );
  AOI21_X2 U152 ( .B1(n304), .B2(n303), .A(n302), .ZN(n309) );
  NAND2_X2 U153 ( .A1(n181), .A2(n97), .ZN(n183) );
  OAI21_X2 U154 ( .B1(n297), .B2(n296), .A(n295), .ZN(n298) );
  AOI21_X2 U155 ( .B1(n210), .B2(n209), .A(n208), .ZN(n211) );
  AOI21_X2 U156 ( .B1(n96), .B2(n202), .A(n201), .ZN(n210) );
  OAI21_X2 U157 ( .B1(b[17]), .B2(a[17]), .A(n99), .ZN(n231) );
  NAND3_X2 U158 ( .A1(n247), .A2(n248), .A3(n115), .ZN(n254) );
  NOR2_X2 U159 ( .A1(n244), .A2(n216), .ZN(n114) );
  NOR2_X2 U160 ( .A1(n269), .A2(n191), .ZN(n123) );
  NAND4_X2 U161 ( .A1(n149), .A2(n148), .A3(n154), .A4(n155), .ZN(n316) );
  AOI21_X2 U162 ( .B1(n157), .B2(n156), .A(n104), .ZN(n158) );
  AOI21_X2 U163 ( .B1(n315), .B2(n147), .A(n317), .ZN(n157) );
  NAND3_X2 U164 ( .A1(n264), .A2(n263), .A3(n262), .ZN(n267) );
  NAND3_X2 U165 ( .A1(n273), .A2(n272), .A3(n271), .ZN(n276) );
  AOI21_X2 U166 ( .B1(n293), .B2(n296), .A(n297), .ZN(n294) );
  AOI21_X2 U167 ( .B1(n313), .B2(n312), .A(n311), .ZN(n314) );
  AND2_X4 U168 ( .A1(n204), .A2(n205), .ZN(n96) );
  XOR2_X2 U169 ( .A(b[10]), .B(a[10]), .Z(n97) );
  XOR2_X2 U170 ( .A(b[9]), .B(a[9]), .Z(n98) );
  XOR2_X2 U171 ( .A(b[18]), .B(a[18]), .Z(n99) );
  XOR2_X2 U172 ( .A(b[29]), .B(a[29]), .Z(n100) );
  AND2_X4 U173 ( .A1(n223), .A2(n225), .ZN(n101) );
  AND2_X4 U174 ( .A1(n147), .A2(n146), .ZN(n102) );
  XOR2_X2 U175 ( .A(b[8]), .B(a[8]), .Z(n103) );
  OAI21_X2 U176 ( .B1(n311), .B2(n312), .A(n100), .ZN(n108) );
  OAI21_X2 U177 ( .B1(n198), .B2(n197), .A(n96), .ZN(n261) );
  AND2_X4 U178 ( .A1(b[31]), .A2(a[31]), .ZN(n104) );
  NAND4_X4 U179 ( .A1(n144), .A2(n143), .A3(n306), .A4(n305), .ZN(n155) );
  NAND4_X4 U180 ( .A1(n186), .A2(n284), .A3(n183), .A4(n285), .ZN(n305) );
  OAI22_X4 U181 ( .A1(n133), .A2(n132), .B1(n162), .B2(n163), .ZN(n166) );
  AOI22_X4 U182 ( .A1(n166), .A2(n134), .B1(b[3]), .B2(a[3]), .ZN(n168) );
  NAND2_X2 U183 ( .A1(b[30]), .A2(a[30]), .ZN(n147) );
  NAND2_X2 U184 ( .A1(b[29]), .A2(a[29]), .ZN(n149) );
  NAND2_X2 U185 ( .A1(b[28]), .A2(a[28]), .ZN(n105) );
  INV_X4 U186 ( .A(n105), .ZN(n311) );
  XNOR2_X2 U187 ( .A(b[28]), .B(a[28]), .ZN(n310) );
  INV_X4 U188 ( .A(n310), .ZN(n312) );
  XNOR2_X2 U189 ( .A(b[27]), .B(a[27]), .ZN(n291) );
  NAND2_X2 U190 ( .A1(b[26]), .A2(a[26]), .ZN(n299) );
  NAND2_X2 U191 ( .A1(b[27]), .A2(a[27]), .ZN(n301) );
  OAI211_X2 U192 ( .C1(n291), .C2(n299), .A(n301), .B(n105), .ZN(n106) );
  NAND2_X2 U193 ( .A1(n143), .A2(n106), .ZN(n148) );
  NAND2_X2 U194 ( .A1(b[25]), .A2(a[25]), .ZN(n300) );
  XNOR2_X2 U195 ( .A(b[26]), .B(a[26]), .ZN(n292) );
  NAND2_X2 U196 ( .A1(n107), .A2(n143), .ZN(n154) );
  XNOR2_X2 U197 ( .A(b[25]), .B(a[25]), .ZN(n289) );
  INV_X4 U198 ( .A(n108), .ZN(n143) );
  XNOR2_X2 U199 ( .A(b[11]), .B(a[11]), .ZN(n187) );
  XNOR2_X2 U200 ( .A(b[24]), .B(a[24]), .ZN(n279) );
  NAND2_X2 U201 ( .A1(b[23]), .A2(a[23]), .ZN(n275) );
  NAND2_X2 U202 ( .A1(b[22]), .A2(a[22]), .ZN(n266) );
  NAND2_X2 U203 ( .A1(b[21]), .A2(a[21]), .ZN(n256) );
  NAND2_X2 U204 ( .A1(b[20]), .A2(a[20]), .ZN(n247) );
  XNOR2_X2 U205 ( .A(b[16]), .B(a[16]), .ZN(n220) );
  XNOR2_X2 U206 ( .A(b[19]), .B(a[19]), .ZN(n230) );
  NAND2_X2 U207 ( .A1(b[18]), .A2(a[18]), .ZN(n232) );
  NAND2_X2 U208 ( .A1(n231), .A2(n232), .ZN(n238) );
  NAND2_X2 U209 ( .A1(b[19]), .A2(a[19]), .ZN(n239) );
  INV_X4 U210 ( .A(n239), .ZN(n109) );
  NAND2_X2 U211 ( .A1(b[16]), .A2(a[16]), .ZN(n223) );
  NAND2_X2 U212 ( .A1(b[17]), .A2(a[17]), .ZN(n225) );
  NAND2_X2 U213 ( .A1(n111), .A2(n238), .ZN(n240) );
  NAND2_X2 U214 ( .A1(n112), .A2(n240), .ZN(n246) );
  XNOR2_X2 U215 ( .A(b[20]), .B(a[20]), .ZN(n244) );
  INV_X4 U216 ( .A(n244), .ZN(n245) );
  NAND2_X2 U217 ( .A1(b[15]), .A2(a[15]), .ZN(n219) );
  NAND3_X2 U218 ( .A1(n219), .A2(n240), .A3(n239), .ZN(n113) );
  XNOR2_X2 U219 ( .A(b[15]), .B(a[15]), .ZN(n216) );
  NAND2_X2 U220 ( .A1(n114), .A2(n246), .ZN(n115) );
  XNOR2_X2 U221 ( .A(b[21]), .B(a[21]), .ZN(n252) );
  INV_X4 U222 ( .A(n252), .ZN(n253) );
  NAND2_X2 U223 ( .A1(b[14]), .A2(a[14]), .ZN(n215) );
  XNOR2_X2 U224 ( .A(b[14]), .B(a[14]), .ZN(n212) );
  NAND2_X2 U225 ( .A1(n117), .A2(n254), .ZN(n118) );
  XNOR2_X2 U226 ( .A(b[22]), .B(a[22]), .ZN(n260) );
  INV_X4 U227 ( .A(n260), .ZN(n263) );
  NAND2_X2 U228 ( .A1(b[13]), .A2(a[13]), .ZN(n207) );
  XNOR2_X2 U229 ( .A(b[13]), .B(a[13]), .ZN(n201) );
  NAND2_X2 U230 ( .A1(n120), .A2(n264), .ZN(n121) );
  NAND3_X2 U231 ( .A1(n266), .A2(n265), .A3(n121), .ZN(n273) );
  XNOR2_X2 U232 ( .A(b[23]), .B(a[23]), .ZN(n269) );
  INV_X4 U233 ( .A(n269), .ZN(n272) );
  NAND2_X2 U234 ( .A1(b[12]), .A2(a[12]), .ZN(n205) );
  NAND3_X2 U235 ( .A1(n273), .A2(n272), .A3(n122), .ZN(n274) );
  XNOR2_X2 U236 ( .A(b[12]), .B(a[12]), .ZN(n191) );
  NAND2_X2 U237 ( .A1(n123), .A2(n273), .ZN(n124) );
  NAND3_X2 U238 ( .A1(n275), .A2(n274), .A3(n124), .ZN(n281) );
  NAND2_X2 U239 ( .A1(b[24]), .A2(a[24]), .ZN(n284) );
  INV_X4 U240 ( .A(n284), .ZN(n125) );
  AOI21_X2 U241 ( .B1(n126), .B2(n281), .A(n125), .ZN(n128) );
  INV_X4 U242 ( .A(n279), .ZN(n280) );
  NAND2_X2 U243 ( .A1(b[11]), .A2(a[11]), .ZN(n193) );
  NAND3_X2 U244 ( .A1(n193), .A2(n274), .A3(n275), .ZN(n127) );
  NAND3_X2 U245 ( .A1(n281), .A2(n280), .A3(n127), .ZN(n285) );
  NAND2_X2 U246 ( .A1(n128), .A2(n285), .ZN(n306) );
  NAND2_X2 U247 ( .A1(b[10]), .A2(a[10]), .ZN(n186) );
  NAND2_X2 U248 ( .A1(b[9]), .A2(a[9]), .ZN(n184) );
  NAND2_X2 U249 ( .A1(b[8]), .A2(a[8]), .ZN(n206) );
  NAND2_X2 U250 ( .A1(b[7]), .A2(a[7]), .ZN(n142) );
  INV_X4 U251 ( .A(a[6]), .ZN(n139) );
  INV_X4 U252 ( .A(b[6]), .ZN(n138) );
  XNOR2_X2 U253 ( .A(b[6]), .B(a[6]), .ZN(n172) );
  INV_X4 U254 ( .A(a[4]), .ZN(n136) );
  INV_X4 U255 ( .A(b[4]), .ZN(n135) );
  XNOR2_X2 U256 ( .A(b[4]), .B(a[4]), .ZN(n167) );
  INV_X4 U257 ( .A(a[2]), .ZN(n133) );
  INV_X4 U258 ( .A(b[2]), .ZN(n132) );
  XNOR2_X2 U259 ( .A(b[2]), .B(a[2]), .ZN(n162) );
  XNOR2_X2 U260 ( .A(b[0]), .B(a[0]), .ZN(n159) );
  INV_X4 U261 ( .A(cin), .ZN(n130) );
  NAND2_X2 U262 ( .A1(b[0]), .A2(a[0]), .ZN(n129) );
  XNOR2_X2 U263 ( .A(b[1]), .B(a[1]), .ZN(n160) );
  INV_X4 U264 ( .A(n160), .ZN(n131) );
  XNOR2_X2 U265 ( .A(b[3]), .B(a[3]), .ZN(n165) );
  INV_X4 U266 ( .A(n165), .ZN(n134) );
  XNOR2_X2 U267 ( .A(b[5]), .B(a[5]), .ZN(n170) );
  INV_X4 U268 ( .A(n170), .ZN(n137) );
  AOI22_X2 U269 ( .A1(n171), .A2(n137), .B1(b[5]), .B2(a[5]), .ZN(n173) );
  OAI22_X2 U270 ( .A1(n139), .A2(n138), .B1(n172), .B2(n173), .ZN(n176) );
  XNOR2_X2 U271 ( .A(b[7]), .B(a[7]), .ZN(n175) );
  INV_X4 U272 ( .A(n175), .ZN(n140) );
  NAND2_X2 U273 ( .A1(n176), .A2(n140), .ZN(n141) );
  NAND2_X2 U274 ( .A1(n142), .A2(n141), .ZN(n177) );
  NAND2_X2 U275 ( .A1(n177), .A2(n103), .ZN(n203) );
  NAND2_X2 U276 ( .A1(n206), .A2(n203), .ZN(n179) );
  NAND2_X2 U277 ( .A1(n179), .A2(n98), .ZN(n197) );
  NAND2_X2 U278 ( .A1(n184), .A2(n197), .ZN(n181) );
  XNOR2_X2 U279 ( .A(b[30]), .B(a[30]), .ZN(n315) );
  INV_X4 U280 ( .A(n315), .ZN(n145) );
  NAND2_X2 U281 ( .A1(n316), .A2(n145), .ZN(n146) );
  XNOR2_X2 U282 ( .A(b[31]), .B(a[31]), .ZN(n317) );
  INV_X4 U283 ( .A(n147), .ZN(n152) );
  INV_X4 U284 ( .A(n148), .ZN(n151) );
  INV_X4 U285 ( .A(n149), .ZN(n150) );
  NAND3_X2 U286 ( .A1(n155), .A2(n154), .A3(n153), .ZN(n156) );
  XOR2_X2 U287 ( .A(n102), .B(n158), .Z(v) );
  XNOR2_X2 U288 ( .A(cin), .B(n159), .ZN(sum[0]) );
  XNOR2_X2 U289 ( .A(n161), .B(n160), .ZN(sum[1]) );
  INV_X4 U290 ( .A(n162), .ZN(n164) );
  XNOR2_X2 U291 ( .A(n164), .B(n163), .ZN(sum[2]) );
  XNOR2_X2 U292 ( .A(n166), .B(n165), .ZN(sum[3]) );
  INV_X4 U293 ( .A(n167), .ZN(n169) );
  XNOR2_X2 U294 ( .A(n169), .B(n168), .ZN(sum[4]) );
  XNOR2_X2 U295 ( .A(n171), .B(n170), .ZN(sum[5]) );
  INV_X4 U296 ( .A(n172), .ZN(n174) );
  XNOR2_X2 U297 ( .A(n174), .B(n173), .ZN(sum[6]) );
  XNOR2_X2 U298 ( .A(n176), .B(n175), .ZN(sum[7]) );
  INV_X4 U299 ( .A(n177), .ZN(n178) );
  XNOR2_X2 U300 ( .A(n103), .B(n178), .ZN(sum[8]) );
  INV_X4 U301 ( .A(n179), .ZN(n180) );
  XNOR2_X2 U302 ( .A(n98), .B(n180), .ZN(sum[9]) );
  INV_X4 U303 ( .A(n181), .ZN(n182) );
  XNOR2_X2 U304 ( .A(n97), .B(n182), .ZN(sum[10]) );
  NAND2_X2 U305 ( .A1(n183), .A2(n186), .ZN(n283) );
  XNOR2_X2 U306 ( .A(n283), .B(n187), .ZN(sum[11]) );
  INV_X4 U307 ( .A(n197), .ZN(n185) );
  NAND2_X2 U308 ( .A1(n184), .A2(n186), .ZN(n192) );
  INV_X4 U309 ( .A(n186), .ZN(n188) );
  INV_X4 U310 ( .A(n187), .ZN(n282) );
  XNOR2_X2 U311 ( .A(n270), .B(n191), .ZN(sum[12]) );
  INV_X4 U312 ( .A(n201), .ZN(n262) );
  NAND2_X2 U313 ( .A1(n190), .A2(n193), .ZN(n200) );
  INV_X4 U314 ( .A(n191), .ZN(n271) );
  NAND2_X2 U315 ( .A1(n200), .A2(n271), .ZN(n198) );
  INV_X4 U316 ( .A(n198), .ZN(n196) );
  INV_X4 U317 ( .A(n192), .ZN(n194) );
  NAND2_X2 U318 ( .A1(n194), .A2(n193), .ZN(n195) );
  NAND2_X2 U319 ( .A1(n196), .A2(n195), .ZN(n204) );
  INV_X4 U320 ( .A(n261), .ZN(n199) );
  XNOR2_X2 U321 ( .A(n262), .B(n199), .ZN(sum[13]) );
  NAND4_X2 U322 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(n209) );
  INV_X4 U323 ( .A(n207), .ZN(n208) );
  INV_X4 U324 ( .A(n211), .ZN(n214) );
  XNOR2_X2 U325 ( .A(n214), .B(n212), .ZN(sum[14]) );
  INV_X4 U326 ( .A(n212), .ZN(n213) );
  NAND2_X2 U327 ( .A1(n214), .A2(n213), .ZN(n257) );
  NAND2_X2 U328 ( .A1(n257), .A2(n215), .ZN(n218) );
  XNOR2_X2 U329 ( .A(n218), .B(n216), .ZN(sum[15]) );
  INV_X4 U330 ( .A(n216), .ZN(n217) );
  NAND2_X2 U331 ( .A1(n218), .A2(n217), .ZN(n249) );
  NAND2_X2 U332 ( .A1(n249), .A2(n219), .ZN(n222) );
  XNOR2_X2 U333 ( .A(n222), .B(n220), .ZN(sum[16]) );
  XNOR2_X2 U334 ( .A(b[17]), .B(a[17]), .ZN(n224) );
  INV_X4 U335 ( .A(n220), .ZN(n221) );
  NAND2_X2 U336 ( .A1(n222), .A2(n221), .ZN(n241) );
  NAND2_X2 U337 ( .A1(n241), .A2(n223), .ZN(n227) );
  XNOR2_X2 U338 ( .A(n224), .B(n227), .ZN(sum[17]) );
  INV_X4 U339 ( .A(n224), .ZN(n228) );
  INV_X4 U340 ( .A(n225), .ZN(n226) );
  AOI21_X2 U341 ( .B1(n228), .B2(n227), .A(n226), .ZN(n229) );
  XNOR2_X2 U342 ( .A(n99), .B(n229), .ZN(sum[18]) );
  INV_X4 U343 ( .A(n230), .ZN(n237) );
  INV_X4 U344 ( .A(n231), .ZN(n235) );
  NAND2_X2 U345 ( .A1(n101), .A2(n241), .ZN(n234) );
  INV_X4 U346 ( .A(n232), .ZN(n233) );
  AOI21_X2 U347 ( .B1(n235), .B2(n234), .A(n233), .ZN(n236) );
  XNOR2_X2 U348 ( .A(n237), .B(n236), .ZN(sum[19]) );
  NAND2_X2 U349 ( .A1(n238), .A2(n237), .ZN(n242) );
  OAI211_X2 U350 ( .C1(n242), .C2(n241), .A(n240), .B(n239), .ZN(n243) );
  XNOR2_X2 U351 ( .A(n244), .B(n243), .ZN(sum[20]) );
  NAND2_X2 U352 ( .A1(n246), .A2(n245), .ZN(n250) );
  OAI211_X2 U353 ( .C1(n250), .C2(n249), .A(n248), .B(n247), .ZN(n251) );
  XNOR2_X2 U354 ( .A(n252), .B(n251), .ZN(sum[21]) );
  NAND2_X2 U355 ( .A1(n254), .A2(n253), .ZN(n258) );
  OAI211_X2 U356 ( .C1(n258), .C2(n257), .A(n256), .B(n255), .ZN(n259) );
  XNOR2_X2 U357 ( .A(n260), .B(n259), .ZN(sum[22]) );
  OAI211_X2 U358 ( .C1(n199), .C2(n267), .A(n266), .B(n265), .ZN(n268) );
  XNOR2_X2 U359 ( .A(n269), .B(n268), .ZN(sum[23]) );
  INV_X4 U360 ( .A(n270), .ZN(n277) );
  OAI211_X2 U361 ( .C1(n277), .C2(n276), .A(n275), .B(n274), .ZN(n278) );
  XNOR2_X2 U362 ( .A(n279), .B(n278), .ZN(sum[24]) );
  NAND2_X2 U363 ( .A1(n281), .A2(n280), .ZN(n287) );
  NAND2_X2 U364 ( .A1(n283), .A2(n282), .ZN(n286) );
  OAI211_X2 U365 ( .C1(n287), .C2(n286), .A(n285), .B(n284), .ZN(n288) );
  XNOR2_X2 U366 ( .A(n289), .B(n288), .ZN(sum[25]) );
  INV_X4 U367 ( .A(n289), .ZN(n307) );
  NAND3_X2 U368 ( .A1(n307), .A2(n306), .A3(n305), .ZN(n290) );
  NAND2_X2 U369 ( .A1(n290), .A2(n300), .ZN(n293) );
  XNOR2_X2 U370 ( .A(n293), .B(n292), .ZN(sum[26]) );
  INV_X4 U371 ( .A(n291), .ZN(n295) );
  INV_X4 U372 ( .A(n292), .ZN(n296) );
  INV_X4 U373 ( .A(n299), .ZN(n297) );
  XNOR2_X2 U374 ( .A(n295), .B(n294), .ZN(sum[27]) );
  INV_X4 U375 ( .A(n298), .ZN(n304) );
  NAND2_X2 U376 ( .A1(n300), .A2(n299), .ZN(n303) );
  INV_X4 U377 ( .A(n301), .ZN(n302) );
  NAND4_X2 U378 ( .A1(n307), .A2(n306), .A3(n305), .A4(n304), .ZN(n308) );
  NAND2_X2 U379 ( .A1(n309), .A2(n308), .ZN(n313) );
  XNOR2_X2 U380 ( .A(n313), .B(n310), .ZN(sum[28]) );
  XNOR2_X2 U381 ( .A(n100), .B(n314), .ZN(sum[29]) );
  XNOR2_X2 U382 ( .A(n316), .B(n315), .ZN(sum[30]) );
  INV_X4 U383 ( .A(n317), .ZN(n318) );
  XNOR2_X2 U384 ( .A(n102), .B(n318), .ZN(sum[31]) );
endmodule

