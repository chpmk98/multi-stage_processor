
module foureach ( x, y, result );
  input [31:0] x;
  input [4:0] y;
  output [35:0] result;
  wire   \ddd/adder[0]/axorb , net81582, net153517, net153524, net153525,
         net153526, net153532, net153533, net153535, net153540, net153541,
         net153543, net153545, net153547, net153548, net153549, net153550,
         net153559, net153560, net153561, net153562, net153598, net153600,
         net153611, net153613, net153617, net153621, net153623, net153630,
         net153633, net153637, net153667, net153669, net153671, net153672,
         net153674, net153696, net153698, net153700, net153701, net153743,
         net153769, net153784, net153788, net153796, net153818, net153823,
         net153828, net153829, net153831, net153832, net153833, net153835,
         net153853, net153856, net153863, net153875, net153876, net153881,
         net153930, net153936, net153937, net153942, net153953, net153958,
         net153959, net153960, net153962, net153967, net153975, net153977,
         net153986, net153996, net154001, net154006, net154025, net154028,
         net154031, net154034, net154038, net154055, net154061, net154083,
         net154091, net154117, net154127, net154143, net154151, net154155,
         net154158, net154166, net154169, net154180, net154205, net154234,
         net154244, net154247, net154250, net154277, net154280, net154283,
         net154285, net154290, net154291, net154293, net154294, net154295,
         net154298, net154308, net154320, net154322, net154323, net154332,
         net154334, net154339, net154341, net154349, net154356, net154391,
         net154423, net154438, net154459, net154462, net154477, net154479,
         net154480, net154481, net154499, net154533, net154534, net154536,
         net154560, net154575, net154578, net154588, net154589, net154595,
         net154602, net154606, net154616, net154619, net154620, net154621,
         net154622, net154623, net154629, net154630, net154642, net154660,
         net154667, net154682, net154685, net154687, net154693, net154694,
         net154696, net154697, net154698, net154699, net154700, net154701,
         net154711, net154719, net154721, net154728, net154731, net154734,
         net154742, net154744, net154760, net154773, net154784, net154786,
         net154788, net154791, net154795, net154796, net154802, net154807,
         net154810, net154815, net154817, net154824, net154826, net154827,
         net154828, net154829, net154842, net154848, net154852, net154855,
         net154856, net154858, net154859, net154861, net154862, net154863,
         net154867, net154877, net154879, net154880, net154885, net154905,
         net154940, net154943, net154947, net154956, net154964, net154968,
         net154971, net155041, net155057, net155112, net155310, net155314,
         net155315, net155324, net155327, net155367, net155379, net155446,
         net155457, net155482, net155484, net155489, net155490, net155493,
         net155496, net155506, net155508, net155511, net155513, net155514,
         net155592, net155624, net155644, net155645, net155657, net155665,
         net155667, net155696, net155697, net155732, net155739, net155744,
         net155773, net155775, net155777, net155780, net155781, net155782,
         net155787, net155791, net155799, net155815, net155819, net155820,
         net155827, net155837, net155835, net155841, net155839, net155859,
         net155857, net155855, net155873, net155869, net155885, net155884,
         net155896, net155985, net156057, net156073, net156089, net156110,
         net156131, net156130, net156156, net156169, net156181, net156180,
         net156333, net156405, net156482, net156541, net156614, net156664,
         net156663, net156708, net156711, net156745, net156760, net156776,
         net156784, net156803, net156811, net156810, net156869, net156989,
         net157038, net157076, net157139, net157159, net157244, net157352,
         net157351, net157350, net157381, net157404, net157416, net157424,
         net157440, net157451, net157450, net157521, net157527, net157532,
         net157531, net157542, net157577, net157576, net157575, net157615,
         net157619, net157644, net157651, net157665, net157664, net157769,
         net157767, net157773, net157836, net157848, net157890, net157892,
         net157939, net158084, net158099, net158117, net158116, net158121,
         net158130, net158146, net158219, net158242, net158256, net158266,
         net158270, net158297, net158305, net158330, net157578, net154033,
         net153968, net154537, net154531, net154529, net154528, net153622,
         net153781, net153778, net153777, net153673, net153631, net154442,
         net154328, net153780, net153779, net154736, net157127, net153952,
         net153951, net156857, net154752, net154745, net156283, net154187,
         net154186, net154179, net154178, net154172, net154171, net154170,
         net157074, net153961, net153699, net156622, net156621, net155865,
         net155863, net154816, net154754, net154753, net154535, net154463,
         net153819, net156462, net155895, net155853, net155851, net155847,
         net154608, net154607, net154530, net154103, net153767, net156806,
         net156805, net156532, net156296, net156148, net156147, net154188,
         net154175, net154094, net154035, net153834, net156047, net154912,
         net154868, net154812, net154811, net154809, net154741, net154460,
         net154911, net154881, net154864, net154814, net153907, net157340,
         net155778, net155735, net155199, net155198, net155039, net154944,
         net154941, net154730, net158324, net157339, net157295, net156537,
         net156533, net154288, net154286, net154276, net154177, net153612,
         net158294, net158293, net158282, net157177, net156792, net156791,
         net156790, net156055, net153697, net153695, net153664, net153663,
         net153662, net153635, net153563, net153551, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918;
  assign result[0] = \ddd/adder[0]/axorb ;
  assign result[34] = net81582;

  NAND2_X2 U649 ( .A1(n2087), .A2(n2086), .ZN(net154620) );
  INV_X8 U650 ( .A(net153996), .ZN(net155985) );
  INV_X4 U651 ( .A(net157339), .ZN(net154286) );
  NAND2_X2 U652 ( .A1(net154701), .A2(net154699), .ZN(n499) );
  NAND3_X2 U653 ( .A1(net156857), .A2(net154682), .A3(n500), .ZN(net154696) );
  INV_X4 U654 ( .A(n499), .ZN(n500) );
  BUF_X4 U655 ( .A(net154700), .Z(net156857) );
  NAND2_X4 U656 ( .A1(n1820), .A2(n1854), .ZN(n1764) );
  XNOR2_X2 U657 ( .A(n1721), .B(n898), .ZN(n501) );
  XNOR2_X2 U658 ( .A(n1865), .B(n503), .ZN(n502) );
  INV_X4 U659 ( .A(n502), .ZN(n1727) );
  INV_X32 U660 ( .A(n1864), .ZN(n503) );
  NOR3_X2 U661 ( .A1(n2037), .A2(n2036), .A3(n2035), .ZN(n2038) );
  NAND2_X2 U662 ( .A1(net154971), .A2(net154968), .ZN(n1906) );
  XNOR2_X2 U663 ( .A(n2272), .B(n504), .ZN(n2275) );
  AND2_X2 U664 ( .A1(n2271), .A2(n2270), .ZN(n504) );
  INV_X8 U665 ( .A(n1703), .ZN(n1749) );
  INV_X2 U666 ( .A(n1413), .ZN(n920) );
  INV_X8 U667 ( .A(n1457), .ZN(n1413) );
  INV_X8 U668 ( .A(n1372), .ZN(n994) );
  XNOR2_X2 U669 ( .A(n585), .B(n505), .ZN(n584) );
  INV_X32 U670 ( .A(n514), .ZN(n505) );
  NAND2_X4 U671 ( .A1(n1289), .A2(n1288), .ZN(n1333) );
  XNOR2_X1 U672 ( .A(n2153), .B(n574), .ZN(result[24]) );
  INV_X2 U673 ( .A(n756), .ZN(n2586) );
  INV_X2 U674 ( .A(net154169), .ZN(n506) );
  NAND2_X2 U675 ( .A1(n2165), .A2(net153533), .ZN(n2185) );
  NAND2_X2 U676 ( .A1(net153937), .A2(net153533), .ZN(n2585) );
  INV_X4 U677 ( .A(n834), .ZN(n507) );
  INV_X4 U678 ( .A(n531), .ZN(n508) );
  INV_X8 U679 ( .A(n531), .ZN(n612) );
  OAI21_X4 U680 ( .B1(n1441), .B2(n1421), .A(n933), .ZN(n1666) );
  AND2_X4 U681 ( .A1(n1404), .A2(n1410), .ZN(n531) );
  NAND2_X4 U682 ( .A1(n1019), .A2(n1020), .ZN(n509) );
  NAND2_X4 U683 ( .A1(n1674), .A2(n1178), .ZN(n540) );
  CLKBUF_X3 U684 ( .A(n1292), .Z(n510) );
  INV_X2 U685 ( .A(n2565), .ZN(n1137) );
  INV_X4 U686 ( .A(n2161), .ZN(n962) );
  INV_X2 U687 ( .A(n2172), .ZN(n1987) );
  NOR2_X1 U688 ( .A1(n2080), .A2(net154711), .ZN(n2041) );
  NAND2_X4 U689 ( .A1(n1395), .A2(n1394), .ZN(n539) );
  NAND2_X2 U690 ( .A1(net154560), .A2(net153968), .ZN(net154760) );
  CLKBUF_X2 U691 ( .A(net154560), .Z(n511) );
  NAND2_X2 U692 ( .A1(n2552), .A2(net156131), .ZN(n2547) );
  NOR2_X4 U693 ( .A1(n1518), .A2(n1517), .ZN(n1520) );
  INV_X4 U694 ( .A(net153961), .ZN(net157074) );
  INV_X8 U695 ( .A(net153699), .ZN(net153961) );
  INV_X4 U696 ( .A(n2842), .ZN(n2843) );
  NAND2_X4 U697 ( .A1(n2842), .A2(n1017), .ZN(n2779) );
  INV_X4 U698 ( .A(n1838), .ZN(n512) );
  INV_X4 U699 ( .A(n512), .ZN(n513) );
  CLKBUF_X2 U700 ( .A(n841), .Z(n514) );
  OAI21_X2 U701 ( .B1(net153535), .B2(n2871), .A(n2873), .ZN(n2887) );
  INV_X1 U702 ( .A(n1502), .ZN(n515) );
  NAND2_X4 U703 ( .A1(n924), .A2(n925), .ZN(n1236) );
  INV_X4 U704 ( .A(net154879), .ZN(net154912) );
  CLKBUF_X3 U705 ( .A(x[7]), .Z(n516) );
  OAI22_X4 U706 ( .A1(n1175), .A2(n2532), .B1(n2704), .B2(net155873), .ZN(n565) );
  INV_X32 U707 ( .A(x[7]), .ZN(net155482) );
  NAND2_X4 U708 ( .A1(n2206), .A2(n2205), .ZN(n1152) );
  INV_X16 U709 ( .A(n2391), .ZN(n2206) );
  OAI21_X4 U710 ( .B1(net154117), .B2(n2457), .A(n2456), .ZN(n2611) );
  AND2_X2 U711 ( .A1(net154968), .A2(net154814), .ZN(n517) );
  NAND2_X4 U712 ( .A1(net154956), .A2(n1118), .ZN(n1001) );
  NAND2_X4 U713 ( .A1(net154956), .A2(n1118), .ZN(n1941) );
  OR2_X2 U714 ( .A1(net154828), .A2(net154964), .ZN(n518) );
  NAND2_X1 U715 ( .A1(n1948), .A2(n1969), .ZN(n519) );
  INV_X8 U716 ( .A(net154685), .ZN(net154699) );
  OAI21_X4 U717 ( .B1(net156462), .B2(net154535), .A(net154734), .ZN(net154685) );
  NAND2_X4 U718 ( .A1(n2828), .A2(n852), .ZN(n2741) );
  NAND2_X4 U719 ( .A1(n2390), .A2(n2389), .ZN(n749) );
  NAND2_X4 U720 ( .A1(n1169), .A2(net153831), .ZN(net154298) );
  NAND2_X4 U721 ( .A1(net154619), .A2(net157836), .ZN(n568) );
  XOR2_X1 U722 ( .A(n830), .B(n2257), .Z(n520) );
  INV_X4 U723 ( .A(n550), .ZN(n551) );
  XNOR2_X2 U724 ( .A(n2323), .B(n2322), .ZN(n2325) );
  NAND2_X4 U725 ( .A1(n2585), .A2(net153936), .ZN(n756) );
  NAND2_X4 U726 ( .A1(n1683), .A2(n1682), .ZN(n538) );
  NOR2_X2 U727 ( .A1(n2575), .A2(n2574), .ZN(n2577) );
  INV_X8 U728 ( .A(net157350), .ZN(net157351) );
  INV_X4 U729 ( .A(n814), .ZN(n815) );
  INV_X4 U730 ( .A(n1704), .ZN(n1707) );
  NAND2_X2 U731 ( .A1(n993), .A2(net157576), .ZN(n523) );
  NAND2_X4 U732 ( .A1(n521), .A2(n522), .ZN(n524) );
  NAND2_X4 U733 ( .A1(n523), .A2(n524), .ZN(n729) );
  INV_X4 U734 ( .A(n993), .ZN(n521) );
  INV_X2 U735 ( .A(net157576), .ZN(n522) );
  INV_X4 U736 ( .A(n729), .ZN(n2139) );
  NAND2_X2 U737 ( .A1(n2287), .A2(n2286), .ZN(n527) );
  NAND2_X4 U738 ( .A1(n525), .A2(n526), .ZN(n528) );
  NAND2_X4 U739 ( .A1(n527), .A2(n528), .ZN(net153967) );
  INV_X4 U740 ( .A(n2287), .ZN(n525) );
  INV_X1 U741 ( .A(n2286), .ZN(n526) );
  INV_X8 U742 ( .A(net153967), .ZN(net154391) );
  INV_X2 U743 ( .A(n2394), .ZN(n820) );
  XNOR2_X1 U744 ( .A(net153524), .B(net153525), .ZN(n2875) );
  NAND2_X2 U745 ( .A1(net156790), .A2(net156791), .ZN(n757) );
  INV_X16 U746 ( .A(n1171), .ZN(n1396) );
  INV_X2 U747 ( .A(n1472), .ZN(n933) );
  NAND2_X4 U748 ( .A1(n2662), .A2(n687), .ZN(n2663) );
  INV_X4 U749 ( .A(n2892), .ZN(n2829) );
  NAND3_X4 U750 ( .A1(net156089), .A2(net153831), .A3(n552), .ZN(n2396) );
  INV_X8 U751 ( .A(n2396), .ZN(n2428) );
  NAND3_X4 U752 ( .A1(n2150), .A2(n2149), .A3(n2148), .ZN(n2142) );
  NAND2_X2 U753 ( .A1(n1165), .A2(n1985), .ZN(net154560) );
  INV_X2 U754 ( .A(net153833), .ZN(n679) );
  XNOR2_X2 U755 ( .A(n569), .B(n1060), .ZN(n853) );
  NAND2_X4 U756 ( .A1(n1040), .A2(n1041), .ZN(n529) );
  BUF_X16 U757 ( .A(n1992), .Z(n825) );
  INV_X4 U758 ( .A(n1668), .ZN(n910) );
  AOI211_X4 U759 ( .C1(n2100), .C2(net157076), .A(n2099), .B(n2098), .ZN(n2101) );
  NAND2_X4 U760 ( .A1(n2666), .A2(net158270), .ZN(n2669) );
  NOR2_X1 U761 ( .A1(net154038), .A2(net156181), .ZN(n2098) );
  NOR2_X4 U762 ( .A1(n2288), .A2(net154391), .ZN(n2292) );
  OAI211_X4 U763 ( .C1(n2518), .C2(n2510), .A(n2511), .B(net153828), .ZN(n2519) );
  INV_X4 U764 ( .A(n1407), .ZN(n1332) );
  NAND2_X1 U765 ( .A1(n1617), .A2(n1736), .ZN(n1541) );
  INV_X8 U766 ( .A(net153828), .ZN(n2631) );
  OAI21_X4 U767 ( .B1(n1223), .B2(n1222), .A(n1221), .ZN(n1258) );
  NAND2_X4 U768 ( .A1(n1011), .A2(n1012), .ZN(n1975) );
  NAND4_X4 U769 ( .A1(n2205), .A2(net154642), .A3(net156169), .A4(net154694), 
        .ZN(n2117) );
  INV_X2 U770 ( .A(n1434), .ZN(n1436) );
  INV_X2 U771 ( .A(n2696), .ZN(n2592) );
  NAND2_X4 U772 ( .A1(n1530), .A2(n1529), .ZN(n1531) );
  INV_X8 U773 ( .A(n1529), .ZN(n1502) );
  NAND2_X4 U774 ( .A1(n1665), .A2(n910), .ZN(n912) );
  XNOR2_X1 U775 ( .A(net154606), .B(net156664), .ZN(n730) );
  NAND2_X2 U776 ( .A1(n1182), .A2(n1939), .ZN(n1940) );
  INV_X8 U777 ( .A(n2477), .ZN(n2702) );
  OAI21_X4 U778 ( .B1(n1966), .B2(n2043), .A(net154693), .ZN(n2287) );
  NAND2_X2 U779 ( .A1(n2855), .A2(n2905), .ZN(n1058) );
  AOI21_X4 U780 ( .B1(n2820), .B2(n2819), .A(n2818), .ZN(n2822) );
  NAND2_X2 U781 ( .A1(n890), .A2(n891), .ZN(n2572) );
  NOR2_X4 U782 ( .A1(n2518), .A2(net156148), .ZN(n552) );
  NAND2_X4 U783 ( .A1(net154616), .A2(net154499), .ZN(n2051) );
  OAI21_X4 U784 ( .B1(n726), .B2(n1408), .A(n1407), .ZN(n1410) );
  NAND3_X1 U785 ( .A1(n686), .A2(net153543), .A3(net153547), .ZN(n2869) );
  NAND2_X2 U786 ( .A1(net154276), .A2(net154277), .ZN(n759) );
  NAND2_X1 U787 ( .A1(n932), .A2(n1666), .ZN(n1668) );
  NAND2_X2 U788 ( .A1(y[3]), .A2(net155791), .ZN(n2705) );
  INV_X4 U789 ( .A(net155837), .ZN(net155827) );
  OAI21_X2 U790 ( .B1(n1601), .B2(n1556), .A(n1555), .ZN(n1557) );
  NAND2_X2 U791 ( .A1(net154629), .A2(n1181), .ZN(n2012) );
  NOR2_X2 U792 ( .A1(x[18]), .A2(net155869), .ZN(n1925) );
  OAI21_X2 U793 ( .B1(n572), .B2(net155857), .A(n1947), .ZN(n1948) );
  INV_X8 U794 ( .A(net153907), .ZN(n771) );
  NOR2_X2 U795 ( .A1(x[26]), .A2(x[25]), .ZN(n2598) );
  OAI21_X1 U796 ( .B1(n2704), .B2(net155839), .A(n2672), .ZN(n2715) );
  OAI21_X1 U797 ( .B1(n1015), .B2(net155827), .A(n1932), .ZN(n2282) );
  OAI21_X1 U798 ( .B1(net155827), .B2(n1427), .A(n1426), .ZN(n1496) );
  NAND2_X2 U799 ( .A1(n639), .A2(n640), .ZN(net154463) );
  INV_X4 U800 ( .A(n630), .ZN(n1299) );
  INV_X16 U801 ( .A(y[0]), .ZN(n632) );
  INV_X16 U802 ( .A(x[6]), .ZN(n631) );
  NAND2_X2 U803 ( .A1(n975), .A2(net157352), .ZN(n977) );
  NAND2_X2 U804 ( .A1(n1788), .A2(n1091), .ZN(n2006) );
  INV_X4 U805 ( .A(n2341), .ZN(n2347) );
  INV_X4 U806 ( .A(net154055), .ZN(n678) );
  INV_X4 U807 ( .A(n2410), .ZN(n2455) );
  INV_X4 U808 ( .A(n2404), .ZN(n2457) );
  INV_X4 U809 ( .A(n2371), .ZN(n917) );
  NAND3_X2 U810 ( .A1(y[1]), .A2(net155739), .A3(x[2]), .ZN(n1217) );
  INV_X4 U811 ( .A(n1582), .ZN(n661) );
  AOI21_X2 U812 ( .B1(n1287), .B2(n1286), .A(n713), .ZN(n1289) );
  NAND3_X2 U813 ( .A1(n1182), .A2(n1926), .A3(n1927), .ZN(n1928) );
  NAND2_X2 U814 ( .A1(n2240), .A2(n2371), .ZN(n2407) );
  NAND2_X2 U815 ( .A1(net157892), .A2(net154943), .ZN(n1050) );
  INV_X4 U816 ( .A(n830), .ZN(n1965) );
  INV_X4 U817 ( .A(net154620), .ZN(net157575) );
  INV_X4 U818 ( .A(n1940), .ZN(n1980) );
  INV_X4 U819 ( .A(n2905), .ZN(n1056) );
  NOR2_X2 U820 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  OAI21_X2 U821 ( .B1(n1346), .B2(n1347), .A(n1363), .ZN(n1674) );
  OAI21_X2 U822 ( .B1(n727), .B2(net155841), .A(n1425), .ZN(n1435) );
  NOR2_X2 U823 ( .A1(n2066), .A2(n2063), .ZN(n2064) );
  OAI21_X2 U824 ( .B1(n733), .B2(net155827), .A(n2249), .ZN(net153986) );
  OAI21_X1 U825 ( .B1(n2414), .B2(net155827), .A(n2413), .ZN(n2571) );
  INV_X4 U826 ( .A(n1366), .ZN(n946) );
  INV_X4 U827 ( .A(n1663), .ZN(n1650) );
  OAI21_X1 U828 ( .B1(n1596), .B2(net155827), .A(n1595), .ZN(n1637) );
  INV_X4 U829 ( .A(n1639), .ZN(n591) );
  OAI21_X1 U830 ( .B1(n829), .B2(net155827), .A(n1722), .ZN(n1864) );
  NAND2_X2 U831 ( .A1(n2302), .A2(n2301), .ZN(n2323) );
  OAI21_X1 U832 ( .B1(net154719), .B2(net155827), .A(n2059), .ZN(n2159) );
  NAND2_X2 U833 ( .A1(n853), .A2(n2830), .ZN(n2753) );
  OAI21_X1 U834 ( .B1(n2804), .B2(net155827), .A(n2803), .ZN(n2907) );
  AOI21_X2 U835 ( .B1(n2901), .B2(n2900), .A(n2899), .ZN(n2906) );
  INV_X4 U836 ( .A(n1316), .ZN(n582) );
  NOR2_X2 U837 ( .A1(n1492), .A2(n1491), .ZN(n1507) );
  CLKBUF_X2 U838 ( .A(net158294), .Z(net158282) );
  INV_X8 U839 ( .A(n771), .ZN(net155873) );
  AND2_X4 U840 ( .A1(x[13]), .A2(net155884), .ZN(n530) );
  INV_X16 U841 ( .A(net155884), .ZN(net155885) );
  BUF_X4 U842 ( .A(n2112), .Z(n900) );
  INV_X4 U843 ( .A(n2705), .ZN(n1183) );
  INV_X2 U844 ( .A(n1617), .ZN(n633) );
  OAI21_X1 U845 ( .B1(net155827), .B2(n2542), .A(n2541), .ZN(net153633) );
  INV_X16 U846 ( .A(x[9]), .ZN(net155496) );
  INV_X16 U847 ( .A(net155847), .ZN(net155841) );
  INV_X4 U848 ( .A(net155837), .ZN(net155835) );
  INV_X4 U849 ( .A(net153637), .ZN(net155837) );
  INV_X2 U850 ( .A(n806), .ZN(n807) );
  INV_X2 U851 ( .A(net154968), .ZN(n738) );
  INV_X4 U852 ( .A(n721), .ZN(n1687) );
  INV_X4 U853 ( .A(n812), .ZN(n2767) );
  INV_X4 U854 ( .A(n804), .ZN(n1039) );
  INV_X4 U855 ( .A(n1169), .ZN(n880) );
  INV_X4 U856 ( .A(n2836), .ZN(n2838) );
  NAND2_X2 U857 ( .A1(n2116), .A2(n2202), .ZN(n2388) );
  INV_X4 U858 ( .A(n2388), .ZN(n2389) );
  INV_X4 U859 ( .A(net154693), .ZN(net156708) );
  INV_X4 U860 ( .A(net154693), .ZN(net154288) );
  AND2_X4 U861 ( .A1(n1276), .A2(n1275), .ZN(n532) );
  INV_X4 U862 ( .A(n2271), .ZN(n619) );
  AND4_X2 U863 ( .A1(net157527), .A2(n568), .A3(n560), .A4(n2074), .ZN(n533)
         );
  AND2_X2 U864 ( .A1(n1736), .A2(n1071), .ZN(n534) );
  AND3_X2 U865 ( .A1(n1781), .A2(n1782), .A3(net155112), .ZN(n535) );
  XNOR2_X2 U866 ( .A(n815), .B(n1656), .ZN(n1665) );
  OAI21_X2 U867 ( .B1(n1996), .B2(n1995), .A(n1994), .ZN(n2417) );
  AND2_X2 U868 ( .A1(n1490), .A2(n1489), .ZN(n536) );
  OR2_X2 U869 ( .A1(x[13]), .A2(x[14]), .ZN(n537) );
  INV_X4 U870 ( .A(n1273), .ZN(n923) );
  OAI211_X2 U871 ( .C1(net154589), .C2(n895), .A(n2000), .B(n2002), .ZN(n2001)
         );
  INV_X4 U872 ( .A(n2001), .ZN(n2252) );
  INV_X4 U873 ( .A(n2781), .ZN(n2709) );
  INV_X8 U874 ( .A(n1004), .ZN(n1411) );
  INV_X4 U875 ( .A(net154339), .ZN(net156156) );
  INV_X4 U876 ( .A(net156156), .ZN(net156869) );
  INV_X4 U877 ( .A(n2609), .ZN(n2613) );
  INV_X8 U878 ( .A(net155853), .ZN(net155851) );
  INV_X8 U879 ( .A(net153767), .ZN(net155853) );
  INV_X4 U880 ( .A(net155869), .ZN(n692) );
  INV_X8 U881 ( .A(net156296), .ZN(net156110) );
  XNOR2_X1 U882 ( .A(n2095), .B(n2325), .ZN(result[23]) );
  NOR2_X2 U883 ( .A1(net153937), .A2(n2174), .ZN(n2176) );
  XNOR2_X1 U884 ( .A(n2378), .B(net153547), .ZN(result[27]) );
  NAND2_X2 U885 ( .A1(n2169), .A2(n2566), .ZN(n1986) );
  NAND2_X4 U886 ( .A1(n1986), .A2(n2284), .ZN(n1960) );
  XNOR2_X2 U887 ( .A(n585), .B(n2286), .ZN(n2319) );
  NOR3_X2 U888 ( .A1(net154760), .A2(n2034), .A3(n2033), .ZN(n2035) );
  NAND2_X2 U889 ( .A1(n2161), .A2(n2160), .ZN(n964) );
  INV_X2 U890 ( .A(n2736), .ZN(n2587) );
  NAND2_X2 U891 ( .A1(n2736), .A2(n549), .ZN(n2328) );
  NAND2_X4 U892 ( .A1(n2327), .A2(n2326), .ZN(n2736) );
  NAND2_X2 U893 ( .A1(n1683), .A2(n1682), .ZN(n2222) );
  NAND2_X4 U894 ( .A1(n1681), .A2(n1740), .ZN(n1682) );
  NAND2_X4 U895 ( .A1(n2023), .A2(n2022), .ZN(n2170) );
  OAI21_X2 U896 ( .B1(n2442), .B2(n2331), .A(n551), .ZN(n2378) );
  OAI22_X4 U897 ( .A1(net155896), .A2(net155592), .B1(net155841), .B2(n1427), 
        .ZN(n1394) );
  INV_X2 U898 ( .A(net154166), .ZN(net154169) );
  INV_X4 U899 ( .A(n695), .ZN(n1963) );
  NAND2_X4 U900 ( .A1(n1877), .A2(n1876), .ZN(n2284) );
  NOR2_X2 U901 ( .A1(n1559), .A2(x[11]), .ZN(n1563) );
  INV_X1 U902 ( .A(n1285), .ZN(n541) );
  INV_X2 U903 ( .A(n541), .ZN(n542) );
  INV_X8 U904 ( .A(n1244), .ZN(n1280) );
  NOR2_X4 U905 ( .A1(n2426), .A2(n2425), .ZN(n2442) );
  OAI21_X2 U906 ( .B1(n2423), .B2(n2442), .A(n2422), .ZN(n2424) );
  NAND2_X2 U907 ( .A1(n1244), .A2(n1283), .ZN(n865) );
  INV_X2 U908 ( .A(n2283), .ZN(n2258) );
  XNOR2_X1 U909 ( .A(n1724), .B(n1727), .ZN(result[14]) );
  OAI21_X2 U910 ( .B1(n2441), .B2(n2442), .A(n2440), .ZN(n2476) );
  NAND2_X4 U911 ( .A1(n2460), .A2(n554), .ZN(n2615) );
  NAND2_X2 U912 ( .A1(net154816), .A2(net154817), .ZN(n639) );
  XNOR2_X2 U913 ( .A(n749), .B(n1021), .ZN(n2509) );
  INV_X1 U914 ( .A(n1857), .ZN(n827) );
  INV_X2 U915 ( .A(n1960), .ZN(n1934) );
  INV_X2 U916 ( .A(n1960), .ZN(n1961) );
  AND2_X4 U917 ( .A1(n1448), .A2(n1447), .ZN(n543) );
  INV_X4 U918 ( .A(n1482), .ZN(n1448) );
  INV_X8 U919 ( .A(n1483), .ZN(n1447) );
  NAND2_X2 U920 ( .A1(n2353), .A2(n519), .ZN(net154283) );
  INV_X4 U921 ( .A(n2768), .ZN(n2770) );
  INV_X4 U922 ( .A(net154817), .ZN(n638) );
  INV_X1 U923 ( .A(n1518), .ZN(n544) );
  XNOR2_X2 U924 ( .A(n1340), .B(n1339), .ZN(n1342) );
  OAI21_X4 U925 ( .B1(n2468), .B2(n2467), .A(n2529), .ZN(n545) );
  NAND2_X4 U926 ( .A1(n1332), .A2(n1331), .ZN(n1335) );
  NOR2_X2 U927 ( .A1(net154031), .A2(n2066), .ZN(n2067) );
  NAND2_X4 U928 ( .A1(n1704), .A2(n1705), .ZN(n546) );
  CLKBUF_X3 U929 ( .A(n1609), .Z(n649) );
  INV_X1 U930 ( .A(n1526), .ZN(n547) );
  INV_X4 U931 ( .A(n547), .ZN(n548) );
  NAND2_X4 U932 ( .A1(net153547), .A2(net153543), .ZN(n2427) );
  BUF_X8 U933 ( .A(n1659), .Z(n1071) );
  XNOR2_X2 U934 ( .A(n2645), .B(n571), .ZN(result[31]) );
  NOR2_X4 U935 ( .A1(n762), .A2(net154177), .ZN(n761) );
  NAND2_X4 U936 ( .A1(n2316), .A2(n2552), .ZN(n549) );
  INV_X2 U937 ( .A(n2545), .ZN(n2316) );
  INV_X2 U938 ( .A(n1571), .ZN(n1421) );
  OAI21_X2 U939 ( .B1(n2110), .B2(n2109), .A(n2108), .ZN(n2153) );
  OAI21_X2 U940 ( .B1(n2110), .B2(n2073), .A(n2072), .ZN(n2095) );
  INV_X2 U941 ( .A(net153540), .ZN(n550) );
  NAND2_X2 U942 ( .A1(n2516), .A2(n2813), .ZN(n2814) );
  INV_X8 U943 ( .A(n1399), .ZN(n660) );
  NAND2_X2 U944 ( .A1(n719), .A2(n716), .ZN(net154856) );
  NAND2_X4 U945 ( .A1(n2189), .A2(n2190), .ZN(n2264) );
  INV_X2 U946 ( .A(net154320), .ZN(net154187) );
  NAND2_X2 U947 ( .A1(n2659), .A2(n2661), .ZN(n2664) );
  AND2_X2 U948 ( .A1(n2429), .A2(n2395), .ZN(n2433) );
  NAND2_X4 U949 ( .A1(n2393), .A2(n2394), .ZN(n2429) );
  INV_X4 U950 ( .A(net154175), .ZN(net154188) );
  INV_X16 U951 ( .A(x[3]), .ZN(net155735) );
  NOR2_X2 U952 ( .A1(x[4]), .A2(x[3]), .ZN(n1443) );
  NAND3_X2 U953 ( .A1(y[1]), .A2(net155739), .A3(x[3]), .ZN(net155732) );
  NAND2_X2 U954 ( .A1(x[0]), .A2(x[3]), .ZN(n1210) );
  INV_X16 U955 ( .A(x[3]), .ZN(net155696) );
  INV_X4 U956 ( .A(x[3]), .ZN(n736) );
  OAI22_X1 U957 ( .A1(net155896), .A2(net155735), .B1(net155841), .B2(
        net155697), .ZN(net155657) );
  OAI21_X2 U958 ( .B1(net155857), .B2(net155697), .A(net155732), .ZN(n1247) );
  NAND2_X2 U959 ( .A1(n1209), .A2(n1444), .ZN(n1198) );
  OAI22_X1 U960 ( .A1(n2705), .A2(net155696), .B1(net155827), .B2(net155697), 
        .ZN(n1352) );
  NAND2_X2 U961 ( .A1(net155696), .A2(net155645), .ZN(n1554) );
  NAND2_X2 U962 ( .A1(net155696), .A2(net155645), .ZN(n558) );
  INV_X4 U963 ( .A(n968), .ZN(n1417) );
  OAI211_X2 U964 ( .C1(n1834), .C2(n835), .A(n1832), .B(net154810), .ZN(n1907)
         );
  CLKBUF_X3 U965 ( .A(net153696), .Z(n553) );
  OAI21_X4 U966 ( .B1(net153598), .B2(n2584), .A(n2878), .ZN(n1022) );
  INV_X4 U967 ( .A(n2403), .ZN(n554) );
  NAND2_X1 U968 ( .A1(n2511), .A2(net154334), .ZN(n698) );
  NAND3_X1 U969 ( .A1(n1168), .A2(net153828), .A3(n687), .ZN(n2513) );
  OAI211_X4 U970 ( .C1(n820), .C2(n2392), .A(n2633), .B(net158270), .ZN(n2526)
         );
  NOR3_X4 U971 ( .A1(n2380), .A2(n2407), .A3(n2379), .ZN(n2382) );
  CLKBUF_X3 U972 ( .A(n1590), .Z(n555) );
  OAI21_X2 U973 ( .B1(n2759), .B2(n2758), .A(n2757), .ZN(n556) );
  INV_X8 U974 ( .A(n751), .ZN(n2758) );
  NAND2_X2 U975 ( .A1(net154619), .A2(net157836), .ZN(n2127) );
  NAND2_X2 U976 ( .A1(n556), .A2(n588), .ZN(n990) );
  INV_X8 U977 ( .A(net158324), .ZN(net156131) );
  INV_X4 U978 ( .A(net158324), .ZN(n617) );
  INV_X1 U979 ( .A(n1307), .ZN(n557) );
  INV_X8 U980 ( .A(net156180), .ZN(net156181) );
  INV_X4 U981 ( .A(n1437), .ZN(n1150) );
  NAND2_X2 U982 ( .A1(n1415), .A2(n1416), .ZN(n1437) );
  INV_X2 U983 ( .A(n2520), .ZN(n2099) );
  NOR2_X2 U984 ( .A1(n816), .A2(n530), .ZN(n930) );
  NAND2_X2 U985 ( .A1(n2357), .A2(n2573), .ZN(n2377) );
  NAND2_X1 U986 ( .A1(n1950), .A2(n1949), .ZN(n666) );
  INV_X2 U987 ( .A(n2043), .ZN(n2134) );
  INV_X4 U988 ( .A(n1093), .ZN(n2465) );
  INV_X16 U989 ( .A(net155865), .ZN(net155863) );
  INV_X1 U990 ( .A(n691), .ZN(n559) );
  NAND2_X2 U991 ( .A1(net154308), .A2(net154280), .ZN(n560) );
  NAND2_X2 U992 ( .A1(net154308), .A2(net154280), .ZN(n561) );
  OAI21_X4 U993 ( .B1(n821), .B2(net155841), .A(n1938), .ZN(net154280) );
  NAND2_X2 U994 ( .A1(net154308), .A2(net154280), .ZN(net154293) );
  NAND2_X4 U995 ( .A1(n1802), .A2(n857), .ZN(n562) );
  BUF_X8 U996 ( .A(n854), .Z(n588) );
  NAND3_X1 U997 ( .A1(net155493), .A2(net155865), .A3(net157351), .ZN(n563) );
  INV_X4 U998 ( .A(n2548), .ZN(n595) );
  NAND2_X2 U999 ( .A1(n605), .A2(net154533), .ZN(n1096) );
  INV_X4 U1000 ( .A(net154499), .ZN(net156333) );
  XNOR2_X2 U1001 ( .A(n1385), .B(n1141), .ZN(n564) );
  XNOR2_X1 U1002 ( .A(n1394), .B(n1411), .ZN(n1385) );
  OAI21_X2 U1003 ( .B1(n1384), .B2(n1383), .A(n823), .ZN(n1141) );
  INV_X2 U1004 ( .A(n1522), .ZN(n1391) );
  INV_X2 U1005 ( .A(n1365), .ZN(n1367) );
  OAI211_X4 U1006 ( .C1(n1834), .C2(n835), .A(n1832), .B(net154810), .ZN(n566)
         );
  INV_X8 U1007 ( .A(net155819), .ZN(n567) );
  INV_X8 U1008 ( .A(net155787), .ZN(net155819) );
  INV_X2 U1009 ( .A(n1649), .ZN(n1616) );
  INV_X8 U1010 ( .A(n2459), .ZN(n2403) );
  NOR2_X2 U1011 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  NAND2_X2 U1012 ( .A1(net157577), .A2(net157578), .ZN(net157836) );
  INV_X4 U1013 ( .A(net156805), .ZN(net156806) );
  NAND2_X1 U1014 ( .A1(n2741), .A2(n2740), .ZN(n569) );
  NAND2_X2 U1015 ( .A1(n2741), .A2(n2740), .ZN(n2742) );
  INV_X2 U1016 ( .A(net154816), .ZN(n637) );
  NAND2_X2 U1017 ( .A1(net154817), .A2(net154816), .ZN(net154535) );
  NOR2_X4 U1018 ( .A1(n1831), .A2(n1888), .ZN(n1832) );
  XOR2_X2 U1019 ( .A(n1647), .B(n721), .Z(n940) );
  INV_X4 U1020 ( .A(net153951), .ZN(net153942) );
  NAND2_X4 U1021 ( .A1(n2336), .A2(n2335), .ZN(n570) );
  NAND2_X2 U1022 ( .A1(n2336), .A2(n2335), .ZN(n2345) );
  XNOR2_X1 U1023 ( .A(n1633), .B(n1649), .ZN(n1635) );
  INV_X4 U1024 ( .A(n935), .ZN(n571) );
  INV_X4 U1025 ( .A(n2749), .ZN(n935) );
  NAND3_X4 U1026 ( .A1(n1369), .A2(n845), .A3(net155859), .ZN(n1322) );
  INV_X8 U1027 ( .A(n844), .ZN(n845) );
  XNOR2_X2 U1028 ( .A(n1001), .B(x[17]), .ZN(n572) );
  INV_X2 U1029 ( .A(net156110), .ZN(n573) );
  INV_X2 U1030 ( .A(n1179), .ZN(n1710) );
  AOI22_X2 U1031 ( .A1(n660), .A2(n1582), .B1(n1580), .B2(n1581), .ZN(n1585)
         );
  INV_X4 U1032 ( .A(n1147), .ZN(n1689) );
  NAND2_X4 U1033 ( .A1(n2721), .A2(n2720), .ZN(n1123) );
  NAND2_X2 U1034 ( .A1(n2721), .A2(n2720), .ZN(n2670) );
  NOR2_X4 U1035 ( .A1(n1472), .A2(n1473), .ZN(n1474) );
  INV_X4 U1036 ( .A(n2305), .ZN(n574) );
  INV_X4 U1037 ( .A(n2324), .ZN(n2305) );
  INV_X2 U1038 ( .A(net153526), .ZN(net153524) );
  OAI211_X2 U1039 ( .C1(n1412), .C2(n673), .A(n612), .B(n1475), .ZN(n575) );
  INV_X8 U1040 ( .A(n1587), .ZN(n1412) );
  NAND2_X2 U1041 ( .A1(n1009), .A2(n1969), .ZN(n1012) );
  NAND2_X2 U1042 ( .A1(n1970), .A2(n1010), .ZN(n1011) );
  NAND2_X4 U1043 ( .A1(n2445), .A2(n2444), .ZN(n576) );
  NAND2_X2 U1044 ( .A1(n1361), .A2(n1360), .ZN(n1364) );
  NOR2_X4 U1045 ( .A1(x[6]), .A2(x[5]), .ZN(n577) );
  NAND2_X4 U1046 ( .A1(n988), .A2(n989), .ZN(n991) );
  NAND2_X1 U1047 ( .A1(n1600), .A2(n1599), .ZN(n578) );
  INV_X1 U1048 ( .A(n2285), .ZN(n579) );
  INV_X4 U1049 ( .A(n579), .ZN(n580) );
  NAND2_X4 U1050 ( .A1(n2510), .A2(n2511), .ZN(n2505) );
  NAND2_X4 U1051 ( .A1(n890), .A2(n891), .ZN(n581) );
  NAND2_X4 U1052 ( .A1(n974), .A2(n674), .ZN(n1180) );
  NOR2_X4 U1053 ( .A1(n558), .A2(n956), .ZN(n974) );
  XNOR2_X2 U1054 ( .A(n582), .B(n1306), .ZN(n1268) );
  INV_X4 U1055 ( .A(n1343), .ZN(n1306) );
  INV_X4 U1056 ( .A(n2479), .ZN(n583) );
  INV_X2 U1057 ( .A(n2345), .ZN(n2346) );
  NAND2_X4 U1058 ( .A1(n1335), .A2(n1334), .ZN(n1336) );
  NAND2_X2 U1059 ( .A1(n798), .A2(n799), .ZN(net153778) );
  INV_X4 U1060 ( .A(net156089), .ZN(net154061) );
  INV_X2 U1061 ( .A(n2501), .ZN(n875) );
  OAI21_X2 U1062 ( .B1(n1966), .B2(n2043), .A(n2524), .ZN(n585) );
  INV_X4 U1063 ( .A(net153550), .ZN(n586) );
  NAND2_X2 U1064 ( .A1(n997), .A2(n998), .ZN(n1000) );
  INV_X1 U1065 ( .A(net156622), .ZN(n609) );
  NAND3_X1 U1066 ( .A1(net154842), .A2(net154560), .A3(net153968), .ZN(n587)
         );
  NAND3_X1 U1067 ( .A1(n1860), .A2(n1859), .A3(n1863), .ZN(n808) );
  INV_X8 U1068 ( .A(n2419), .ZN(n937) );
  INV_X2 U1069 ( .A(n1770), .ZN(n1683) );
  XNOR2_X2 U1070 ( .A(n1890), .B(n1720), .ZN(n1885) );
  OAI21_X2 U1071 ( .B1(n1817), .B2(net155841), .A(n1760), .ZN(n1891) );
  OAI22_X1 U1072 ( .A1(n2705), .A2(n1818), .B1(n1817), .B2(net155827), .ZN(
        n1823) );
  XNOR2_X2 U1073 ( .A(net154328), .B(net153829), .ZN(n589) );
  INV_X16 U1074 ( .A(net156148), .ZN(net153829) );
  NAND2_X1 U1075 ( .A1(net154824), .A2(net156622), .ZN(n610) );
  OAI22_X4 U1076 ( .A1(net155896), .A2(n2362), .B1(net155841), .B2(n2472), 
        .ZN(n2444) );
  INV_X2 U1077 ( .A(n707), .ZN(n706) );
  NAND2_X4 U1078 ( .A1(n1769), .A2(n1768), .ZN(n1740) );
  NAND2_X4 U1079 ( .A1(net156784), .A2(n2289), .ZN(n2291) );
  XOR2_X2 U1080 ( .A(n2405), .B(n2406), .Z(n590) );
  OAI22_X4 U1081 ( .A1(net155885), .A2(n2362), .B1(net155855), .B2(n2472), 
        .ZN(n2406) );
  XNOR2_X2 U1082 ( .A(n591), .B(n1638), .ZN(n1644) );
  NOR2_X4 U1083 ( .A1(x[10]), .A2(x[9]), .ZN(n592) );
  NOR2_X4 U1084 ( .A1(x[10]), .A2(x[9]), .ZN(n593) );
  NAND3_X2 U1085 ( .A1(net158305), .A2(n2516), .A3(net157527), .ZN(n1082) );
  NAND4_X2 U1086 ( .A1(n744), .A2(n1839), .A3(n745), .A4(n746), .ZN(n594) );
  OAI211_X2 U1087 ( .C1(n2066), .C2(net158146), .A(n2523), .B(net157527), .ZN(
        n855) );
  INV_X4 U1088 ( .A(n2815), .ZN(n2816) );
  OAI22_X2 U1089 ( .A1(n2158), .A2(n2314), .B1(n2157), .B2(n2301), .ZN(n2161)
         );
  INV_X8 U1090 ( .A(n1376), .ZN(n1582) );
  INV_X8 U1091 ( .A(n2236), .ZN(n2194) );
  OAI21_X4 U1092 ( .B1(n1016), .B2(n2193), .A(n2192), .ZN(n2236) );
  INV_X4 U1093 ( .A(net154811), .ZN(net154741) );
  INV_X4 U1094 ( .A(net154033), .ZN(net156805) );
  OAI211_X2 U1095 ( .C1(n801), .C2(n2027), .A(n2026), .B(n2172), .ZN(n2029) );
  OAI21_X2 U1096 ( .B1(n801), .B2(n1825), .A(n2026), .ZN(n1851) );
  INV_X4 U1097 ( .A(n2167), .ZN(n596) );
  INV_X4 U1098 ( .A(n2319), .ZN(n2167) );
  INV_X1 U1099 ( .A(n1228), .ZN(n597) );
  INV_X2 U1100 ( .A(n597), .ZN(n598) );
  NAND2_X4 U1101 ( .A1(n1748), .A2(n837), .ZN(n1752) );
  NAND2_X2 U1102 ( .A1(net154941), .A2(net155513), .ZN(net155644) );
  INV_X4 U1103 ( .A(n895), .ZN(n599) );
  INV_X4 U1104 ( .A(n2417), .ZN(n895) );
  INV_X1 U1105 ( .A(net154828), .ZN(n600) );
  INV_X8 U1106 ( .A(net154810), .ZN(net154828) );
  NAND2_X4 U1107 ( .A1(n2418), .A2(n599), .ZN(n601) );
  NAND2_X2 U1108 ( .A1(n2418), .A2(n599), .ZN(n2515) );
  BUF_X32 U1109 ( .A(n1497), .Z(n602) );
  OAI21_X4 U1110 ( .B1(n836), .B2(net155855), .A(n1328), .ZN(n1303) );
  NAND2_X4 U1111 ( .A1(x[5]), .A2(net155884), .ZN(n1328) );
  INV_X1 U1112 ( .A(n1363), .ZN(n603) );
  XNOR2_X2 U1113 ( .A(net154911), .B(net154912), .ZN(n604) );
  INV_X1 U1114 ( .A(n1736), .ZN(n1737) );
  NAND2_X4 U1115 ( .A1(net154807), .A2(n781), .ZN(n605) );
  INV_X8 U1116 ( .A(n1303), .ZN(n1331) );
  INV_X8 U1117 ( .A(n1906), .ZN(n1910) );
  INV_X8 U1118 ( .A(n1170), .ZN(n606) );
  NAND3_X4 U1119 ( .A1(net153829), .A2(n908), .A3(net153831), .ZN(n2666) );
  INV_X8 U1120 ( .A(n1177), .ZN(n1178) );
  CLKBUF_X3 U1121 ( .A(net157381), .Z(n607) );
  NAND2_X1 U1122 ( .A1(net154809), .A2(net154700), .ZN(net154867) );
  NAND2_X2 U1123 ( .A1(n2163), .A2(n2162), .ZN(n2164) );
  INV_X8 U1124 ( .A(n1350), .ZN(n1363) );
  INV_X2 U1125 ( .A(n1000), .ZN(n624) );
  NAND2_X2 U1126 ( .A1(n623), .A2(n624), .ZN(n626) );
  NAND2_X4 U1127 ( .A1(n608), .A2(n609), .ZN(n611) );
  NAND2_X4 U1128 ( .A1(n610), .A2(n611), .ZN(net154536) );
  INV_X4 U1129 ( .A(net154824), .ZN(n608) );
  INV_X2 U1130 ( .A(net154536), .ZN(net154528) );
  NAND3_X2 U1131 ( .A1(net154827), .A2(net154682), .A3(n600), .ZN(n1977) );
  NAND2_X4 U1132 ( .A1(n1216), .A2(n1217), .ZN(n1224) );
  OAI22_X4 U1133 ( .A1(n1175), .A2(n2089), .B1(n2250), .B2(net155869), .ZN(
        n2114) );
  XNOR2_X2 U1134 ( .A(n1527), .B(n1525), .ZN(n1390) );
  NAND2_X4 U1135 ( .A1(n1701), .A2(n1702), .ZN(n1802) );
  NAND2_X2 U1136 ( .A1(n2260), .A2(n2259), .ZN(n702) );
  INV_X4 U1137 ( .A(n2775), .ZN(n1076) );
  INV_X1 U1138 ( .A(net153563), .ZN(net158293) );
  NAND2_X4 U1139 ( .A1(n2712), .A2(n2711), .ZN(n2713) );
  NAND2_X2 U1140 ( .A1(n791), .A2(net154298), .ZN(n788) );
  INV_X2 U1141 ( .A(net154158), .ZN(net154155) );
  NAND2_X4 U1142 ( .A1(n1134), .A2(n1794), .ZN(n851) );
  BUF_X8 U1143 ( .A(n1723), .Z(n829) );
  NAND2_X2 U1144 ( .A1(n2198), .A2(n2197), .ZN(n615) );
  NAND2_X4 U1145 ( .A1(n613), .A2(n614), .ZN(n616) );
  NAND2_X4 U1146 ( .A1(n615), .A2(n616), .ZN(n2391) );
  INV_X4 U1147 ( .A(n2198), .ZN(n613) );
  INV_X2 U1148 ( .A(n2197), .ZN(n614) );
  OAI21_X4 U1149 ( .B1(n1016), .B2(n2125), .A(n2124), .ZN(n2197) );
  CLKBUF_X2 U1150 ( .A(n2391), .Z(n1176) );
  INV_X2 U1151 ( .A(n2443), .ZN(n1067) );
  INV_X2 U1152 ( .A(n606), .ZN(n889) );
  OAI21_X4 U1153 ( .B1(n812), .B2(net153853), .A(n2764), .ZN(n2648) );
  INV_X8 U1154 ( .A(n2648), .ZN(n2849) );
  NAND2_X4 U1155 ( .A1(n1069), .A2(n1070), .ZN(n2445) );
  NAND2_X2 U1156 ( .A1(n2718), .A2(n2717), .ZN(n2719) );
  INV_X8 U1157 ( .A(n1172), .ZN(n1175) );
  INV_X8 U1158 ( .A(n1172), .ZN(n1174) );
  NAND4_X2 U1159 ( .A1(n2887), .A2(n2886), .A3(n2884), .A4(n2885), .ZN(n2888)
         );
  NAND2_X4 U1160 ( .A1(y[1]), .A2(n770), .ZN(net155820) );
  NAND2_X2 U1161 ( .A1(n2014), .A2(n2271), .ZN(n620) );
  NAND2_X4 U1162 ( .A1(n618), .A2(n619), .ZN(n621) );
  NAND2_X4 U1163 ( .A1(n620), .A2(n621), .ZN(n2032) );
  INV_X4 U1164 ( .A(n2014), .ZN(n618) );
  NAND2_X2 U1165 ( .A1(n2268), .A2(n2269), .ZN(n2014) );
  INV_X4 U1166 ( .A(n2032), .ZN(n2288) );
  NOR2_X2 U1167 ( .A1(net154588), .A2(net156482), .ZN(n790) );
  NAND2_X4 U1168 ( .A1(net154685), .A2(net154694), .ZN(n2244) );
  INV_X4 U1169 ( .A(net157773), .ZN(n622) );
  INV_X8 U1170 ( .A(net155985), .ZN(net157773) );
  NOR2_X2 U1171 ( .A1(n1865), .A2(n1864), .ZN(n1866) );
  NAND2_X4 U1172 ( .A1(n949), .A2(net155506), .ZN(n1483) );
  CLKBUF_X3 U1173 ( .A(n2074), .Z(n969) );
  NAND2_X1 U1174 ( .A1(n1290), .A2(n1000), .ZN(n625) );
  NAND2_X2 U1175 ( .A1(n625), .A2(n626), .ZN(n737) );
  INV_X1 U1176 ( .A(n1290), .ZN(n623) );
  OAI21_X4 U1177 ( .B1(n2382), .B2(n2381), .A(n2409), .ZN(n2383) );
  INV_X2 U1178 ( .A(net153743), .ZN(net157038) );
  INV_X4 U1179 ( .A(n1418), .ZN(n1113) );
  NAND2_X4 U1180 ( .A1(n754), .A2(net158121), .ZN(n753) );
  INV_X8 U1181 ( .A(n2746), .ZN(n2747) );
  NAND2_X2 U1182 ( .A1(net154175), .A2(n2517), .ZN(net154179) );
  OAI21_X4 U1183 ( .B1(n1708), .B2(net155644), .A(x[6]), .ZN(n1369) );
  NAND2_X2 U1184 ( .A1(n1369), .A2(n845), .ZN(n1427) );
  NAND2_X4 U1185 ( .A1(n2664), .A2(n2663), .ZN(net153832) );
  INV_X2 U1186 ( .A(n1334), .ZN(n1293) );
  NAND2_X4 U1187 ( .A1(n1377), .A2(n1405), .ZN(n1334) );
  NAND2_X4 U1188 ( .A1(n694), .A2(n1755), .ZN(n1847) );
  INV_X4 U1189 ( .A(n2499), .ZN(n2500) );
  AOI22_X4 U1190 ( .A1(n1382), .A2(n1326), .B1(n1382), .B2(net155869), .ZN(
        n1409) );
  BUF_X16 U1191 ( .A(n1404), .Z(n823) );
  NOR2_X4 U1192 ( .A1(n1747), .A2(n530), .ZN(n627) );
  INV_X8 U1193 ( .A(n1745), .ZN(n1747) );
  NOR2_X4 U1194 ( .A1(n2431), .A2(n2482), .ZN(n2432) );
  INV_X8 U1195 ( .A(n1422), .ZN(n1472) );
  NAND2_X4 U1196 ( .A1(n982), .A2(n983), .ZN(n1583) );
  INV_X2 U1197 ( .A(n2484), .ZN(n2485) );
  NAND2_X2 U1198 ( .A1(n2188), .A2(n883), .ZN(n2189) );
  INV_X4 U1199 ( .A(n699), .ZN(n2897) );
  INV_X4 U1200 ( .A(n2848), .ZN(n2766) );
  NAND2_X2 U1201 ( .A1(n2616), .A2(n2501), .ZN(n877) );
  INV_X1 U1202 ( .A(n2723), .ZN(n2639) );
  NAND3_X1 U1203 ( .A1(n552), .A2(net153831), .A3(net156089), .ZN(n2446) );
  OAI21_X1 U1204 ( .B1(n1503), .B2(n1502), .A(n507), .ZN(n628) );
  XNOR2_X2 U1205 ( .A(n1203), .B(n1202), .ZN(n629) );
  OAI211_X4 U1206 ( .C1(net155624), .C2(n631), .A(y[1]), .B(n632), .ZN(n630)
         );
  NAND2_X1 U1207 ( .A1(n1617), .A2(n1505), .ZN(n635) );
  NAND2_X2 U1208 ( .A1(n633), .A2(n634), .ZN(n636) );
  NAND2_X2 U1209 ( .A1(n635), .A2(n636), .ZN(n1458) );
  INV_X4 U1210 ( .A(n1505), .ZN(n634) );
  OAI22_X1 U1211 ( .A1(n2705), .A2(net155482), .B1(n727), .B2(net155827), .ZN(
        n1505) );
  NAND3_X4 U1212 ( .A1(n1494), .A2(n1678), .A3(n1493), .ZN(n1177) );
  NAND2_X2 U1213 ( .A1(n637), .A2(n638), .ZN(n640) );
  AOI22_X4 U1214 ( .A1(n1991), .A2(n2222), .B1(n2218), .B2(n2074), .ZN(n2253)
         );
  NOR2_X2 U1215 ( .A1(n1049), .A2(n863), .ZN(n1991) );
  OR2_X2 U1216 ( .A1(n2735), .A2(n2734), .ZN(n641) );
  NAND2_X2 U1217 ( .A1(n641), .A2(n2733), .ZN(n2759) );
  INV_X4 U1218 ( .A(n1835), .ZN(n1099) );
  NAND3_X2 U1219 ( .A1(n808), .A2(n2026), .A3(n1862), .ZN(n919) );
  NAND2_X4 U1220 ( .A1(n1824), .A2(n1823), .ZN(n2026) );
  INV_X32 U1221 ( .A(x[1]), .ZN(n748) );
  INV_X1 U1222 ( .A(n1397), .ZN(n1401) );
  NAND2_X4 U1223 ( .A1(n865), .A2(n866), .ZN(n1310) );
  NAND3_X2 U1224 ( .A1(n1304), .A2(n1294), .A3(net155859), .ZN(n1243) );
  NAND2_X1 U1225 ( .A1(n2616), .A2(n2614), .ZN(n2622) );
  INV_X4 U1226 ( .A(n605), .ZN(net156663) );
  INV_X4 U1227 ( .A(net154460), .ZN(n642) );
  INV_X8 U1228 ( .A(net154460), .ZN(net158297) );
  INV_X8 U1229 ( .A(net153612), .ZN(net154276) );
  NAND2_X4 U1230 ( .A1(n2489), .A2(n2488), .ZN(n2490) );
  INV_X4 U1231 ( .A(n2411), .ZN(n2443) );
  XNOR2_X2 U1232 ( .A(net154905), .B(n644), .ZN(n643) );
  XOR2_X2 U1233 ( .A(net154280), .B(net156537), .Z(n644) );
  INV_X1 U1234 ( .A(net153962), .ZN(net153958) );
  NAND3_X2 U1235 ( .A1(n2517), .A2(n687), .A3(n2510), .ZN(n2512) );
  NAND2_X2 U1236 ( .A1(n2377), .A2(n2576), .ZN(n647) );
  NAND2_X4 U1237 ( .A1(n645), .A2(n646), .ZN(n648) );
  NAND2_X4 U1238 ( .A1(n647), .A2(n648), .ZN(net153547) );
  INV_X4 U1239 ( .A(n2377), .ZN(n645) );
  INV_X1 U1240 ( .A(n2576), .ZN(n646) );
  INV_X4 U1241 ( .A(net153547), .ZN(net153548) );
  NAND2_X2 U1242 ( .A1(n1127), .A2(net156614), .ZN(n976) );
  INV_X1 U1243 ( .A(net156614), .ZN(net157352) );
  INV_X8 U1244 ( .A(net156462), .ZN(net156169) );
  NAND2_X4 U1245 ( .A1(n1549), .A2(n1553), .ZN(n1037) );
  NAND2_X4 U1246 ( .A1(n2203), .A2(n2206), .ZN(n650) );
  NAND3_X4 U1247 ( .A1(n2204), .A2(n2234), .A3(n651), .ZN(n2408) );
  INV_X4 U1248 ( .A(n650), .ZN(n651) );
  OAI22_X1 U1249 ( .A1(n567), .A2(net155835), .B1(n2705), .B2(net155775), .ZN(
        n1275) );
  NAND3_X1 U1250 ( .A1(net155775), .A2(net157450), .A3(net156745), .ZN(n1708)
         );
  NAND2_X2 U1251 ( .A1(n563), .A2(net155489), .ZN(n654) );
  NAND2_X4 U1252 ( .A1(n652), .A2(n653), .ZN(n655) );
  NAND2_X4 U1253 ( .A1(n654), .A2(n655), .ZN(n1456) );
  INV_X4 U1254 ( .A(net155490), .ZN(n652) );
  INV_X4 U1255 ( .A(net155489), .ZN(n653) );
  NAND2_X4 U1256 ( .A1(n1660), .A2(n1736), .ZN(n959) );
  NAND2_X4 U1257 ( .A1(n952), .A2(n953), .ZN(n955) );
  NAND2_X4 U1258 ( .A1(n818), .A2(net153856), .ZN(n2655) );
  NAND2_X2 U1259 ( .A1(n2808), .A2(n576), .ZN(n2504) );
  INV_X8 U1260 ( .A(n1804), .ZN(n835) );
  CLKBUF_X3 U1261 ( .A(n826), .Z(n656) );
  INV_X2 U1262 ( .A(net154602), .ZN(net156803) );
  NAND2_X2 U1263 ( .A1(n2139), .A2(net154602), .ZN(n2137) );
  INV_X32 U1264 ( .A(x[4]), .ZN(n735) );
  NAND2_X2 U1265 ( .A1(n2199), .A2(n2202), .ZN(n2234) );
  CLKBUF_X2 U1266 ( .A(n2199), .Z(n1003) );
  NAND2_X2 U1267 ( .A1(n1357), .A2(n1356), .ZN(n1523) );
  XNOR2_X2 U1268 ( .A(n1356), .B(n1171), .ZN(n1348) );
  NAND2_X1 U1269 ( .A1(n1617), .A2(n1459), .ZN(n658) );
  NAND2_X2 U1270 ( .A1(n633), .A2(n657), .ZN(n659) );
  NAND2_X2 U1271 ( .A1(n658), .A2(n659), .ZN(n1506) );
  INV_X1 U1272 ( .A(n1459), .ZN(n657) );
  NAND2_X4 U1273 ( .A1(n1504), .A2(n1660), .ZN(n1459) );
  NAND3_X2 U1274 ( .A1(n2753), .A2(n2751), .A3(net153669), .ZN(n2756) );
  NAND2_X4 U1275 ( .A1(net155506), .A2(n949), .ZN(n918) );
  NAND2_X1 U1276 ( .A1(n859), .A2(net154143), .ZN(n2867) );
  OAI211_X1 U1277 ( .C1(n2070), .C2(n2043), .A(n560), .B(n2042), .ZN(n2044) );
  AND3_X2 U1278 ( .A1(n2872), .A2(net153533), .A3(net153532), .ZN(n2874) );
  NAND3_X4 U1279 ( .A1(n2097), .A2(net156760), .A3(n1087), .ZN(n2082) );
  NAND2_X4 U1280 ( .A1(n2309), .A2(n2308), .ZN(n2326) );
  INV_X4 U1281 ( .A(n2210), .ZN(n2333) );
  NAND3_X4 U1282 ( .A1(n1213), .A2(net155327), .A3(net155777), .ZN(n1200) );
  INV_X4 U1283 ( .A(n1192), .ZN(n1223) );
  NAND2_X2 U1284 ( .A1(n1399), .A2(n1582), .ZN(n662) );
  NAND2_X4 U1285 ( .A1(n660), .A2(n661), .ZN(n663) );
  NAND2_X4 U1286 ( .A1(n663), .A2(n662), .ZN(n1004) );
  NAND2_X4 U1287 ( .A1(n664), .A2(n665), .ZN(n667) );
  NAND2_X4 U1288 ( .A1(n666), .A2(n667), .ZN(net156784) );
  INV_X2 U1289 ( .A(n1950), .ZN(n664) );
  INV_X1 U1290 ( .A(n1949), .ZN(n665) );
  INV_X8 U1291 ( .A(net156784), .ZN(net153968) );
  XOR2_X1 U1292 ( .A(n1355), .B(n1171), .Z(n1357) );
  NAND2_X1 U1293 ( .A1(n2694), .A2(n2693), .ZN(n670) );
  NAND2_X4 U1294 ( .A1(n668), .A2(n669), .ZN(n671) );
  NAND2_X4 U1295 ( .A1(n670), .A2(n671), .ZN(n2746) );
  INV_X2 U1296 ( .A(n2694), .ZN(n668) );
  INV_X4 U1297 ( .A(n2693), .ZN(n669) );
  INV_X1 U1298 ( .A(n1080), .ZN(n2693) );
  INV_X4 U1299 ( .A(n2627), .ZN(n1166) );
  NAND3_X2 U1300 ( .A1(n747), .A2(n748), .A3(n714), .ZN(n672) );
  INV_X8 U1301 ( .A(x[2]), .ZN(n747) );
  INV_X4 U1302 ( .A(n1588), .ZN(n673) );
  XNOR2_X1 U1303 ( .A(n1694), .B(n1566), .ZN(n721) );
  NAND2_X4 U1304 ( .A1(n756), .A2(net153532), .ZN(net153697) );
  INV_X8 U1305 ( .A(n1167), .ZN(n2649) );
  NOR4_X4 U1306 ( .A1(x[6]), .A2(x[5]), .A3(x[8]), .A4(x[7]), .ZN(n674) );
  INV_X4 U1307 ( .A(n1748), .ZN(n1889) );
  INV_X8 U1308 ( .A(net153560), .ZN(net153562) );
  NAND2_X4 U1309 ( .A1(net154341), .A2(n969), .ZN(n2016) );
  NAND2_X2 U1310 ( .A1(net154642), .A2(net154616), .ZN(n675) );
  NAND2_X4 U1311 ( .A1(n676), .A2(n2118), .ZN(net154807) );
  INV_X4 U1312 ( .A(n675), .ZN(n676) );
  INV_X8 U1313 ( .A(net155327), .ZN(net155379) );
  INV_X16 U1314 ( .A(net157890), .ZN(net154943) );
  BUF_X4 U1315 ( .A(n1885), .Z(n898) );
  INV_X1 U1316 ( .A(n2844), .ZN(n677) );
  OAI21_X2 U1317 ( .B1(n1473), .B2(n932), .A(n1807), .ZN(n1468) );
  NAND3_X4 U1318 ( .A1(net154642), .A2(net154694), .A3(net156169), .ZN(n2128)
         );
  NAND3_X4 U1319 ( .A1(n1755), .A2(n771), .A3(n694), .ZN(n1716) );
  NAND2_X1 U1320 ( .A1(n516), .A2(net153769), .ZN(n1425) );
  NAND2_X4 U1321 ( .A1(net155884), .A2(n516), .ZN(n1398) );
  NAND2_X4 U1322 ( .A1(x[8]), .A2(x[7]), .ZN(n1371) );
  NAND2_X2 U1323 ( .A1(n841), .A2(net154602), .ZN(n2186) );
  NOR2_X2 U1324 ( .A1(n1259), .A2(n1258), .ZN(n1260) );
  INV_X4 U1325 ( .A(net153622), .ZN(net158116) );
  INV_X4 U1326 ( .A(net154537), .ZN(net154619) );
  XNOR2_X2 U1327 ( .A(n678), .B(net154250), .ZN(n773) );
  INV_X4 U1328 ( .A(net154205), .ZN(net154250) );
  NAND3_X1 U1329 ( .A1(net155775), .A2(net157451), .A3(net157440), .ZN(
        net155457) );
  NOR2_X2 U1330 ( .A1(net154188), .A2(net158330), .ZN(net154186) );
  NAND2_X4 U1331 ( .A1(n2847), .A2(n2846), .ZN(n2854) );
  NOR2_X4 U1332 ( .A1(n1569), .A2(n839), .ZN(n1570) );
  NAND2_X2 U1333 ( .A1(n2156), .A2(n2329), .ZN(n2158) );
  INV_X4 U1334 ( .A(n2507), .ZN(n2394) );
  INV_X2 U1335 ( .A(n939), .ZN(n680) );
  INV_X4 U1336 ( .A(n939), .ZN(n1079) );
  OAI21_X4 U1337 ( .B1(n2185), .B2(n2184), .A(n2183), .ZN(n2213) );
  XNOR2_X1 U1338 ( .A(n1315), .B(n1343), .ZN(n1317) );
  INV_X2 U1339 ( .A(n1226), .ZN(n1201) );
  NAND2_X1 U1340 ( .A1(n1226), .A2(n1288), .ZN(n1222) );
  NAND3_X1 U1341 ( .A1(n1220), .A2(n1288), .A3(n1226), .ZN(n1221) );
  NAND3_X2 U1342 ( .A1(n1405), .A2(n1403), .A3(n1377), .ZN(n1378) );
  NAND2_X4 U1343 ( .A1(n2514), .A2(n937), .ZN(n938) );
  NAND2_X4 U1344 ( .A1(n1758), .A2(n1145), .ZN(n1100) );
  INV_X4 U1345 ( .A(n1911), .ZN(n1815) );
  NAND2_X4 U1346 ( .A1(n911), .A2(n912), .ZN(n1672) );
  NAND2_X2 U1347 ( .A1(n849), .A2(n1285), .ZN(n1279) );
  NAND3_X1 U1348 ( .A1(n595), .A2(n2517), .A3(n687), .ZN(n2630) );
  XNOR2_X2 U1349 ( .A(n827), .B(n1855), .ZN(n2024) );
  INV_X4 U1350 ( .A(net158121), .ZN(net153559) );
  OAI21_X1 U1351 ( .B1(n2176), .B2(n2175), .A(n574), .ZN(n2182) );
  NAND2_X4 U1352 ( .A1(n1353), .A2(n1352), .ZN(n1516) );
  INV_X4 U1353 ( .A(n1224), .ZN(n996) );
  NAND2_X2 U1354 ( .A1(n2084), .A2(n2083), .ZN(n683) );
  NAND2_X4 U1355 ( .A1(n681), .A2(n682), .ZN(n684) );
  NAND2_X4 U1356 ( .A1(n683), .A2(n684), .ZN(net154462) );
  INV_X4 U1357 ( .A(n2083), .ZN(n681) );
  INV_X4 U1358 ( .A(n2084), .ZN(n682) );
  NAND3_X2 U1359 ( .A1(net154462), .A2(n2239), .A3(n2202), .ZN(n2203) );
  INV_X16 U1360 ( .A(net154462), .ZN(net154694) );
  OAI22_X2 U1361 ( .A1(net155896), .A2(net155624), .B1(n1148), .B2(net155841), 
        .ZN(n1366) );
  XNOR2_X1 U1362 ( .A(n2076), .B(net157532), .ZN(n685) );
  NAND2_X4 U1363 ( .A1(net154697), .A2(net154696), .ZN(n2076) );
  NAND2_X2 U1364 ( .A1(n685), .A2(net154623), .ZN(n2520) );
  INV_X8 U1365 ( .A(net154694), .ZN(net157531) );
  OAI21_X4 U1366 ( .B1(net154288), .B2(net157139), .A(net154290), .ZN(
        net158219) );
  NAND2_X4 U1367 ( .A1(x[17]), .A2(n1947), .ZN(n1918) );
  NAND2_X4 U1368 ( .A1(x[17]), .A2(n1915), .ZN(n1947) );
  OAI21_X4 U1369 ( .B1(net155839), .B2(n2093), .A(n2058), .ZN(net154623) );
  NAND2_X4 U1370 ( .A1(net155379), .A2(n943), .ZN(n1294) );
  OAI21_X1 U1371 ( .B1(n2540), .B2(n2539), .A(n2538), .ZN(n819) );
  NOR2_X2 U1372 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  NAND2_X4 U1373 ( .A1(n581), .A2(n2571), .ZN(n686) );
  AOI21_X4 U1374 ( .B1(n2866), .B2(n2865), .A(n2864), .ZN(n2870) );
  NAND2_X4 U1375 ( .A1(n529), .A2(n2386), .ZN(n687) );
  INV_X1 U1376 ( .A(n1475), .ZN(n688) );
  NAND2_X4 U1377 ( .A1(n689), .A2(n690), .ZN(n1836) );
  INV_X4 U1378 ( .A(n1937), .ZN(n691) );
  INV_X1 U1379 ( .A(n1175), .ZN(n693) );
  NAND2_X4 U1380 ( .A1(n691), .A2(n692), .ZN(n689) );
  NAND2_X1 U1381 ( .A1(x[16]), .A2(n693), .ZN(n690) );
  NAND2_X2 U1382 ( .A1(n2367), .A2(n2366), .ZN(n2409) );
  NAND2_X2 U1383 ( .A1(n2642), .A2(net156541), .ZN(n2812) );
  INV_X4 U1384 ( .A(n1808), .ZN(n856) );
  NAND2_X2 U1385 ( .A1(n1695), .A2(n847), .ZN(n1684) );
  NAND2_X2 U1386 ( .A1(n1715), .A2(n704), .ZN(n694) );
  OAI21_X4 U1387 ( .B1(net156283), .B2(net155869), .A(net154880), .ZN(n772) );
  INV_X2 U1388 ( .A(n1837), .ZN(n970) );
  NAND2_X2 U1389 ( .A1(n1959), .A2(n1958), .ZN(n695) );
  NAND3_X2 U1390 ( .A1(n760), .A2(net154171), .A3(net154172), .ZN(n696) );
  OAI21_X4 U1391 ( .B1(n2314), .B2(n2102), .A(n2101), .ZN(net154660) );
  NAND2_X2 U1392 ( .A1(n2315), .A2(n1169), .ZN(n881) );
  NAND3_X2 U1393 ( .A1(n887), .A2(n1281), .A3(n943), .ZN(n697) );
  OAI22_X4 U1394 ( .A1(net155896), .A2(n1839), .B1(n1015), .B2(net155841), 
        .ZN(n1902) );
  XNOR2_X2 U1395 ( .A(n2713), .B(n2782), .ZN(n699) );
  OAI21_X1 U1396 ( .B1(n2804), .B2(net155841), .A(n2706), .ZN(n2908) );
  NAND2_X2 U1397 ( .A1(net154534), .A2(net154536), .ZN(n2521) );
  NAND2_X4 U1398 ( .A1(net154536), .A2(net154534), .ZN(n2065) );
  NAND2_X4 U1399 ( .A1(net154308), .A2(net154280), .ZN(n2524) );
  NOR2_X4 U1400 ( .A1(n1413), .A2(net155857), .ZN(n1414) );
  INV_X16 U1401 ( .A(net155859), .ZN(net155857) );
  INV_X4 U1402 ( .A(n2789), .ZN(n2895) );
  INV_X4 U1403 ( .A(n1612), .ZN(n984) );
  INV_X4 U1404 ( .A(n711), .ZN(n1610) );
  NOR2_X4 U1405 ( .A1(n2122), .A2(n2600), .ZN(n2123) );
  NAND2_X4 U1406 ( .A1(n2121), .A2(n2120), .ZN(n2600) );
  INV_X4 U1407 ( .A(n2399), .ZN(n2400) );
  OAI21_X4 U1408 ( .B1(net154288), .B2(net157139), .A(net154290), .ZN(
        net153612) );
  NAND2_X2 U1409 ( .A1(n813), .A2(n1220), .ZN(n1194) );
  NAND2_X4 U1410 ( .A1(n1454), .A2(n1455), .ZN(net157350) );
  NAND2_X2 U1411 ( .A1(net154094), .A2(net154175), .ZN(net156532) );
  NOR2_X4 U1412 ( .A1(n1258), .A2(n1259), .ZN(n700) );
  INV_X4 U1413 ( .A(n700), .ZN(n1225) );
  INV_X4 U1414 ( .A(n2761), .ZN(n2266) );
  NAND2_X2 U1415 ( .A1(n2262), .A2(n2261), .ZN(n701) );
  NOR2_X4 U1416 ( .A1(n701), .A2(n702), .ZN(n703) );
  NAND2_X4 U1417 ( .A1(n2257), .A2(n1165), .ZN(n2260) );
  NOR2_X4 U1418 ( .A1(x[13]), .A2(x[14]), .ZN(n704) );
  NOR3_X4 U1419 ( .A1(n2747), .A2(n2834), .A3(n2748), .ZN(n705) );
  INV_X1 U1420 ( .A(n1741), .ZN(n707) );
  NAND2_X4 U1421 ( .A1(n962), .A2(n963), .ZN(n965) );
  AOI21_X4 U1422 ( .B1(n734), .B2(net155847), .A(n709), .ZN(n708) );
  INV_X4 U1423 ( .A(n708), .ZN(n2386) );
  AND2_X2 U1424 ( .A1(x[23]), .A2(net153769), .ZN(n709) );
  INV_X1 U1425 ( .A(n2250), .ZN(n734) );
  INV_X8 U1426 ( .A(net155847), .ZN(net155839) );
  NAND4_X2 U1427 ( .A1(n2259), .A2(n2261), .A3(n2260), .A4(n2262), .ZN(n710)
         );
  INV_X1 U1428 ( .A(n2902), .ZN(n2903) );
  NAND2_X4 U1429 ( .A1(n2802), .A2(n2911), .ZN(n2902) );
  INV_X2 U1430 ( .A(n1002), .ZN(n2225) );
  OAI21_X4 U1431 ( .B1(net155855), .B2(n1763), .A(n1607), .ZN(n711) );
  INV_X4 U1432 ( .A(n1610), .ZN(n712) );
  AOI21_X4 U1433 ( .B1(net155863), .B2(n1184), .A(n714), .ZN(n713) );
  INV_X4 U1434 ( .A(n713), .ZN(n1189) );
  INV_X32 U1435 ( .A(x[0]), .ZN(n714) );
  NAND2_X4 U1436 ( .A1(y[1]), .A2(net155739), .ZN(n1184) );
  NAND3_X4 U1437 ( .A1(net153701), .A2(n2762), .A3(n1103), .ZN(net153698) );
  NAND2_X4 U1438 ( .A1(n1231), .A2(n999), .ZN(n1265) );
  OAI22_X4 U1439 ( .A1(n1175), .A2(n2089), .B1(n2250), .B2(net155869), .ZN(
        n715) );
  INV_X8 U1440 ( .A(n2088), .ZN(n2250) );
  INV_X8 U1441 ( .A(n1586), .ZN(n1692) );
  INV_X8 U1442 ( .A(net154028), .ZN(net154025) );
  NOR2_X4 U1443 ( .A1(n1978), .A2(net154858), .ZN(n716) );
  AND2_X2 U1444 ( .A1(n717), .A2(net154728), .ZN(n718) );
  INV_X4 U1445 ( .A(net154859), .ZN(n717) );
  AND2_X4 U1446 ( .A1(n717), .A2(net154863), .ZN(n719) );
  NOR2_X2 U1447 ( .A1(n1978), .A2(n720), .ZN(net154731) );
  NAND2_X1 U1448 ( .A1(n717), .A2(n767), .ZN(n720) );
  INV_X8 U1449 ( .A(net154858), .ZN(n767) );
  NAND3_X4 U1450 ( .A1(net155310), .A2(net154861), .A3(net154862), .ZN(n1978)
         );
  NAND2_X4 U1451 ( .A1(n1977), .A2(n1976), .ZN(n1999) );
  BUF_X8 U1452 ( .A(n994), .Z(n1151) );
  INV_X2 U1453 ( .A(net153623), .ZN(net153617) );
  NOR2_X4 U1454 ( .A1(n2880), .A2(net153517), .ZN(n2881) );
  NAND2_X2 U1455 ( .A1(n2543), .A2(net153743), .ZN(n1031) );
  INV_X4 U1456 ( .A(n2543), .ZN(n1030) );
  NAND2_X1 U1457 ( .A1(n2406), .A2(n2405), .ZN(n2456) );
  OAI21_X4 U1458 ( .B1(n900), .B2(net155839), .A(n2090), .ZN(n2140) );
  INV_X4 U1459 ( .A(n722), .ZN(net154816) );
  NOR2_X4 U1460 ( .A1(net154864), .A2(net155855), .ZN(n723) );
  NOR2_X1 U1461 ( .A1(net155885), .A2(net154863), .ZN(n724) );
  NOR2_X4 U1462 ( .A1(n723), .A2(n724), .ZN(n722) );
  INV_X8 U1463 ( .A(net154881), .ZN(net154864) );
  XNOR2_X2 U1464 ( .A(net154170), .B(net156089), .ZN(n725) );
  NAND2_X4 U1465 ( .A1(n725), .A2(net153953), .ZN(net153951) );
  AOI22_X4 U1466 ( .A1(n1326), .A2(n1382), .B1(n1382), .B2(net155869), .ZN(
        n726) );
  INV_X1 U1467 ( .A(n728), .ZN(n727) );
  INV_X1 U1468 ( .A(n1326), .ZN(n728) );
  OAI22_X1 U1469 ( .A1(n2705), .A2(net155484), .B1(net155827), .B2(n1461), 
        .ZN(n1510) );
  NAND2_X2 U1470 ( .A1(n1151), .A2(n920), .ZN(n1461) );
  INV_X4 U1471 ( .A(net153545), .ZN(net153780) );
  INV_X2 U1472 ( .A(n2266), .ZN(n1103) );
  INV_X8 U1473 ( .A(net154463), .ZN(net156621) );
  NAND2_X4 U1474 ( .A1(n1754), .A2(n1753), .ZN(n1758) );
  XNOR2_X1 U1475 ( .A(n2205), .B(n2091), .ZN(net154621) );
  OAI22_X4 U1476 ( .A1(net155885), .A2(n2089), .B1(n2250), .B2(net155855), 
        .ZN(n2198) );
  NAND2_X4 U1477 ( .A1(n732), .A2(n2197), .ZN(n2240) );
  BUF_X8 U1478 ( .A(net156462), .Z(net157244) );
  INV_X8 U1479 ( .A(n2005), .ZN(n1790) );
  NAND2_X4 U1480 ( .A1(n882), .A2(n881), .ZN(n2545) );
  NOR2_X4 U1481 ( .A1(x[7]), .A2(x[8]), .ZN(n731) );
  NOR3_X2 U1482 ( .A1(n1840), .A2(x[9]), .A3(n957), .ZN(n1449) );
  NAND3_X1 U1483 ( .A1(net155775), .A2(net155773), .A3(net157440), .ZN(n957)
         );
  AND4_X4 U1484 ( .A1(n2043), .A2(n568), .A3(n617), .A4(n561), .ZN(n2138) );
  INV_X8 U1485 ( .A(n1829), .ZN(n1895) );
  INV_X8 U1486 ( .A(net154698), .ZN(net154499) );
  OAI22_X2 U1487 ( .A1(net155885), .A2(n2089), .B1(n2250), .B2(net155855), 
        .ZN(n732) );
  INV_X1 U1488 ( .A(n734), .ZN(n733) );
  OAI21_X4 U1489 ( .B1(n567), .B2(net155863), .A(net155799), .ZN(net155815) );
  NAND4_X4 U1490 ( .A1(n735), .A2(n736), .A3(net155041), .A4(y[2]), .ZN(n1560)
         );
  NOR2_X4 U1491 ( .A1(x[19]), .A2(x[20]), .ZN(net154728) );
  INV_X4 U1492 ( .A(n737), .ZN(n1203) );
  NAND3_X2 U1493 ( .A1(n943), .A2(n1281), .A3(n1923), .ZN(n2004) );
  INV_X4 U1494 ( .A(n1117), .ZN(n1281) );
  NAND2_X4 U1495 ( .A1(n1715), .A2(n704), .ZN(n1776) );
  NOR2_X4 U1496 ( .A1(n1901), .A2(n738), .ZN(n739) );
  INV_X4 U1497 ( .A(n739), .ZN(n1140) );
  NOR2_X4 U1498 ( .A1(x[17]), .A2(x[18]), .ZN(n765) );
  NAND2_X4 U1499 ( .A1(n955), .A2(n954), .ZN(n2834) );
  NAND2_X4 U1500 ( .A1(n2849), .A2(n2848), .ZN(n2828) );
  NAND3_X2 U1501 ( .A1(n1099), .A2(n1753), .A3(n1754), .ZN(n1101) );
  NAND2_X4 U1502 ( .A1(n1127), .A2(n1126), .ZN(n1129) );
  INV_X1 U1503 ( .A(n1816), .ZN(n1126) );
  OAI21_X4 U1504 ( .B1(n2266), .B2(n919), .A(net153696), .ZN(n2320) );
  NAND2_X2 U1505 ( .A1(net154629), .A2(net154630), .ZN(n1182) );
  NOR2_X4 U1506 ( .A1(n546), .A2(n1610), .ZN(n740) );
  INV_X4 U1507 ( .A(n740), .ZN(n893) );
  NOR2_X4 U1508 ( .A1(n741), .A2(n708), .ZN(net156482) );
  INV_X2 U1509 ( .A(n2387), .ZN(n741) );
  NAND2_X4 U1510 ( .A1(n1111), .A2(n2581), .ZN(n2729) );
  NAND2_X2 U1511 ( .A1(n2570), .A2(n1124), .ZN(n742) );
  INV_X4 U1512 ( .A(n742), .ZN(n1098) );
  XNOR2_X2 U1513 ( .A(n961), .B(n886), .ZN(n743) );
  INV_X8 U1514 ( .A(n743), .ZN(net153831) );
  NAND2_X4 U1515 ( .A1(n589), .A2(net153986), .ZN(net153540) );
  NAND3_X2 U1516 ( .A1(n2807), .A2(n2808), .A3(net158266), .ZN(n2768) );
  NAND4_X4 U1517 ( .A1(n744), .A2(n1839), .A3(n745), .A4(n746), .ZN(n2005) );
  INV_X4 U1518 ( .A(x[16]), .ZN(n744) );
  INV_X4 U1519 ( .A(x[10]), .ZN(n745) );
  INV_X32 U1520 ( .A(x[9]), .ZN(n746) );
  OAI21_X4 U1521 ( .B1(n2682), .B2(n2683), .A(n2681), .ZN(n2716) );
  INV_X2 U1522 ( .A(n2785), .ZN(n2682) );
  OAI21_X4 U1523 ( .B1(net154294), .B2(net154295), .A(n2351), .ZN(n2575) );
  INV_X2 U1524 ( .A(net158099), .ZN(net154294) );
  OAI22_X2 U1525 ( .A1(net155484), .A2(net154103), .B1(n1461), .B2(net153767), 
        .ZN(n1464) );
  NAND2_X4 U1526 ( .A1(n2656), .A2(n2657), .ZN(n2890) );
  NAND4_X2 U1527 ( .A1(n2709), .A2(n2783), .A3(n2784), .A4(n2785), .ZN(n2712)
         );
  NAND2_X4 U1528 ( .A1(n1815), .A2(n1814), .ZN(n1967) );
  XNOR2_X2 U1529 ( .A(net154247), .B(n784), .ZN(net153875) );
  OAI22_X2 U1530 ( .A1(net155775), .A2(net154103), .B1(net155787), .B2(
        net153767), .ZN(n1230) );
  NAND3_X4 U1531 ( .A1(n747), .A2(n748), .A3(n714), .ZN(net155314) );
  XNOR2_X2 U1532 ( .A(n2405), .B(n2406), .ZN(net154117) );
  NAND3_X2 U1533 ( .A1(n1336), .A2(n1403), .A3(n1337), .ZN(n1338) );
  NAND2_X4 U1534 ( .A1(n972), .A2(net157381), .ZN(net155057) );
  NAND2_X4 U1535 ( .A1(n1584), .A2(n1585), .ZN(n1586) );
  OAI21_X4 U1536 ( .B1(n2570), .B2(n750), .A(n1124), .ZN(n751) );
  INV_X4 U1537 ( .A(n2737), .ZN(n750) );
  INV_X4 U1538 ( .A(n2738), .ZN(n1124) );
  NOR2_X4 U1539 ( .A1(n1117), .A2(n1042), .ZN(n1784) );
  OAI21_X4 U1540 ( .B1(net154864), .B2(net153907), .A(net154880), .ZN(
        net154911) );
  NAND2_X2 U1541 ( .A1(net156792), .A2(n757), .ZN(net81582) );
  INV_X1 U1542 ( .A(net158294), .ZN(net156791) );
  INV_X2 U1543 ( .A(net158293), .ZN(net158294) );
  INV_X4 U1544 ( .A(net153635), .ZN(net156790) );
  NAND2_X1 U1545 ( .A1(net153635), .A2(net158282), .ZN(net156792) );
  XNOR2_X2 U1546 ( .A(net153525), .B(net153526), .ZN(net153563) );
  NOR2_X2 U1547 ( .A1(net153562), .A2(net153563), .ZN(net153561) );
  OAI21_X4 U1548 ( .B1(net153662), .B2(net153663), .A(net153664), .ZN(
        net153635) );
  OAI21_X4 U1549 ( .B1(n753), .B2(n752), .A(net153667), .ZN(net153664) );
  NOR2_X4 U1550 ( .A1(n758), .A2(n755), .ZN(n752) );
  INV_X4 U1551 ( .A(net153672), .ZN(n755) );
  INV_X4 U1552 ( .A(net153796), .ZN(n758) );
  INV_X4 U1553 ( .A(net153669), .ZN(n754) );
  NAND2_X2 U1554 ( .A1(net156055), .A2(net153667), .ZN(net153663) );
  OR2_X2 U1555 ( .A1(net153673), .A2(net153674), .ZN(net156055) );
  NOR4_X2 U1556 ( .A1(net157177), .A2(net153695), .A3(net153673), .A4(
        net153551), .ZN(net153662) );
  INV_X4 U1557 ( .A(net153696), .ZN(net153551) );
  NOR2_X4 U1558 ( .A1(net153550), .A2(net153551), .ZN(net153549) );
  INV_X4 U1559 ( .A(net153697), .ZN(net153695) );
  INV_X2 U1560 ( .A(net153695), .ZN(net157159) );
  INV_X8 U1561 ( .A(net154349), .ZN(net153937) );
  AOI21_X2 U1562 ( .B1(net157074), .B2(net153698), .A(net153700), .ZN(
        net157177) );
  NAND2_X4 U1563 ( .A1(net156533), .A2(n764), .ZN(n760) );
  NAND3_X2 U1564 ( .A1(n760), .A2(net154171), .A3(net154172), .ZN(net154170)
         );
  INV_X4 U1565 ( .A(n763), .ZN(n764) );
  NAND2_X4 U1566 ( .A1(n761), .A2(n759), .ZN(n763) );
  NAND2_X4 U1567 ( .A1(net154276), .A2(net154277), .ZN(net158305) );
  INV_X8 U1568 ( .A(n643), .ZN(net157139) );
  BUF_X8 U1569 ( .A(net154286), .Z(net156537) );
  XNOR2_X2 U1570 ( .A(net154283), .B(net156537), .ZN(net154885) );
  NAND3_X4 U1571 ( .A1(net154815), .A2(net154286), .A3(net154868), .ZN(
        net154700) );
  INV_X1 U1572 ( .A(net156537), .ZN(net156989) );
  NAND3_X1 U1573 ( .A1(net154814), .A2(net154815), .A3(net154286), .ZN(
        net154826) );
  XNOR2_X2 U1574 ( .A(net154911), .B(net154879), .ZN(net157339) );
  NAND2_X2 U1575 ( .A1(net157527), .A2(n2517), .ZN(net154177) );
  INV_X4 U1576 ( .A(net154588), .ZN(net157295) );
  INV_X8 U1577 ( .A(net156131), .ZN(net154588) );
  INV_X8 U1578 ( .A(net153613), .ZN(net158324) );
  INV_X4 U1579 ( .A(net154180), .ZN(n762) );
  NOR2_X2 U1580 ( .A1(net154179), .A2(n762), .ZN(net154178) );
  INV_X4 U1581 ( .A(net156532), .ZN(net156533) );
  NAND2_X4 U1582 ( .A1(net154630), .A2(net154629), .ZN(n766) );
  XNOR2_X2 U1583 ( .A(n766), .B(net154863), .ZN(net154881) );
  INV_X16 U1584 ( .A(net154944), .ZN(net154629) );
  NAND3_X4 U1585 ( .A1(n767), .A2(n768), .A3(n765), .ZN(net154944) );
  NAND2_X2 U1586 ( .A1(n765), .A2(net154728), .ZN(net154802) );
  NOR3_X4 U1587 ( .A1(net157424), .A2(x[12]), .A3(x[11]), .ZN(n768) );
  INV_X8 U1588 ( .A(net154730), .ZN(net154630) );
  NAND3_X2 U1589 ( .A1(net154941), .A2(net155199), .A3(net157340), .ZN(
        net154730) );
  NOR4_X4 U1590 ( .A1(x[6]), .A2(x[5]), .A3(x[8]), .A4(x[7]), .ZN(net157340)
         );
  INV_X8 U1591 ( .A(net155039), .ZN(net155199) );
  NAND2_X4 U1592 ( .A1(net157892), .A2(net155199), .ZN(net155367) );
  NAND3_X4 U1593 ( .A1(net155775), .A2(net155773), .A3(net156745), .ZN(
        net155039) );
  NAND3_X4 U1594 ( .A1(net155775), .A2(net155773), .A3(net157665), .ZN(
        net157890) );
  INV_X32 U1595 ( .A(x[2]), .ZN(net155773) );
  INV_X32 U1596 ( .A(x[1]), .ZN(net155775) );
  INV_X8 U1597 ( .A(net155778), .ZN(net154941) );
  NAND4_X4 U1598 ( .A1(net154943), .A2(net154941), .A3(n1553), .A4(n731), .ZN(
        net154855) );
  NAND2_X4 U1599 ( .A1(net155379), .A2(net154941), .ZN(net155667) );
  NAND2_X4 U1600 ( .A1(net155735), .A2(net155198), .ZN(net155778) );
  INV_X16 U1601 ( .A(x[4]), .ZN(net155198) );
  NAND2_X4 U1602 ( .A1(net155735), .A2(net155645), .ZN(net157404) );
  NAND2_X4 U1603 ( .A1(net154947), .A2(net154940), .ZN(net154859) );
  NAND2_X4 U1604 ( .A1(net154814), .A2(n604), .ZN(n769) );
  OAI21_X4 U1605 ( .B1(net154812), .B2(n769), .A(net154809), .ZN(net154811) );
  INV_X8 U1606 ( .A(net155057), .ZN(net154814) );
  CLKBUF_X3 U1607 ( .A(net154814), .Z(net156614) );
  INV_X32 U1608 ( .A(n771), .ZN(net155869) );
  NAND2_X4 U1609 ( .A1(y[1]), .A2(n770), .ZN(net153907) );
  INV_X32 U1610 ( .A(y[0]), .ZN(n770) );
  BUF_X8 U1611 ( .A(net154864), .Z(net156283) );
  XNOR2_X1 U1612 ( .A(net156057), .B(net154863), .ZN(net154788) );
  NAND2_X4 U1613 ( .A1(net154741), .A2(net154700), .ZN(net154460) );
  NAND2_X4 U1614 ( .A1(net154741), .A2(net154700), .ZN(net154616) );
  INV_X4 U1615 ( .A(net154815), .ZN(net154812) );
  NAND3_X2 U1616 ( .A1(net154285), .A2(net157381), .A3(net154877), .ZN(
        net154868) );
  NAND2_X4 U1617 ( .A1(n772), .A2(net156047), .ZN(net154809) );
  NAND2_X4 U1618 ( .A1(net154809), .A2(net154810), .ZN(net154745) );
  INV_X1 U1619 ( .A(net154912), .ZN(net156047) );
  NOR2_X4 U1620 ( .A1(net154320), .A2(net154188), .ZN(net158099) );
  NAND3_X2 U1621 ( .A1(net156806), .A2(net153622), .A3(net156110), .ZN(
        net154094) );
  NAND3_X2 U1622 ( .A1(net158305), .A2(net157527), .A3(net154094), .ZN(
        net154127) );
  NAND2_X4 U1623 ( .A1(net153623), .A2(net154094), .ZN(net154295) );
  NAND3_X2 U1624 ( .A1(net154158), .A2(net154178), .A3(net154094), .ZN(
        net154172) );
  NAND3_X2 U1625 ( .A1(net154034), .A2(net156806), .A3(net156110), .ZN(
        net153611) );
  NAND3_X4 U1626 ( .A1(net153622), .A2(net156806), .A3(net156110), .ZN(
        net153996) );
  INV_X8 U1627 ( .A(net154035), .ZN(net156296) );
  NAND2_X2 U1628 ( .A1(net154660), .A2(n573), .ZN(net157769) );
  NOR4_X2 U1629 ( .A1(net154031), .A2(net154025), .A3(net156181), .A4(
        net156296), .ZN(net154595) );
  NAND2_X4 U1630 ( .A1(net157578), .A2(net157577), .ZN(net154035) );
  NAND2_X4 U1631 ( .A1(net156811), .A2(net153829), .ZN(net154175) );
  INV_X16 U1632 ( .A(net156147), .ZN(net156148) );
  NOR2_X4 U1633 ( .A1(net154298), .A2(net156148), .ZN(net158330) );
  NOR3_X4 U1634 ( .A1(net153832), .A2(net153833), .A3(net156148), .ZN(
        net153823) );
  INV_X4 U1635 ( .A(net153834), .ZN(net156147) );
  XNOR2_X2 U1636 ( .A(net154442), .B(n773), .ZN(net153834) );
  NAND2_X4 U1637 ( .A1(net154607), .A2(net154608), .ZN(net154530) );
  BUF_X8 U1638 ( .A(net154530), .Z(net156760) );
  INV_X1 U1639 ( .A(net154530), .ZN(net154711) );
  OAI211_X4 U1640 ( .C1(net154528), .C2(net154529), .A(net154530), .B(
        net154537), .ZN(net153622) );
  XNOR2_X2 U1641 ( .A(net154752), .B(net156169), .ZN(net154607) );
  NAND2_X4 U1642 ( .A1(n778), .A2(n779), .ZN(net156462) );
  NAND2_X4 U1643 ( .A1(n776), .A2(n777), .ZN(n779) );
  INV_X8 U1644 ( .A(net154736), .ZN(n777) );
  INV_X1 U1645 ( .A(n777), .ZN(net158130) );
  INV_X4 U1646 ( .A(net154791), .ZN(n776) );
  NAND2_X2 U1647 ( .A1(net154791), .A2(net154736), .ZN(n778) );
  OAI21_X4 U1648 ( .B1(net154719), .B2(net155841), .A(n774), .ZN(net154608) );
  NAND2_X4 U1649 ( .A1(net157939), .A2(net154608), .ZN(net154038) );
  INV_X4 U1650 ( .A(net154608), .ZN(net154786) );
  NAND2_X2 U1651 ( .A1(x[19]), .A2(net153769), .ZN(n774) );
  INV_X16 U1652 ( .A(net155896), .ZN(net153769) );
  INV_X32 U1653 ( .A(net155895), .ZN(net155896) );
  INV_X32 U1654 ( .A(net154103), .ZN(net155895) );
  NAND2_X4 U1655 ( .A1(y[2]), .A2(n775), .ZN(net154103) );
  INV_X4 U1656 ( .A(y[3]), .ZN(n775) );
  NAND2_X2 U1657 ( .A1(y[4]), .A2(n775), .ZN(net153637) );
  INV_X16 U1658 ( .A(net155851), .ZN(net155847) );
  NAND2_X4 U1659 ( .A1(y[3]), .A2(net155739), .ZN(net153767) );
  INV_X32 U1660 ( .A(y[2]), .ZN(net155739) );
  OAI21_X4 U1661 ( .B1(net158297), .B2(net156622), .A(n781), .ZN(net154754) );
  OAI21_X4 U1662 ( .B1(net154753), .B2(net154745), .A(net154754), .ZN(
        net154752) );
  INV_X8 U1663 ( .A(n780), .ZN(n781) );
  NAND2_X4 U1664 ( .A1(net154807), .A2(n781), .ZN(net154606) );
  NAND3_X2 U1665 ( .A1(n2046), .A2(net156857), .A3(n781), .ZN(net154753) );
  NAND2_X2 U1666 ( .A1(net154534), .A2(n781), .ZN(net154531) );
  INV_X4 U1667 ( .A(net154535), .ZN(n780) );
  INV_X16 U1668 ( .A(net156621), .ZN(net156622) );
  INV_X16 U1669 ( .A(net156622), .ZN(net154642) );
  NOR3_X2 U1670 ( .A1(net157244), .A2(net157531), .A3(net156622), .ZN(
        net154459) );
  NAND2_X4 U1671 ( .A1(net156621), .A2(net156169), .ZN(net154698) );
  OAI21_X4 U1672 ( .B1(net158297), .B2(net156333), .A(net157644), .ZN(
        net154697) );
  INV_X32 U1673 ( .A(net155859), .ZN(net155855) );
  INV_X32 U1674 ( .A(net155863), .ZN(net155859) );
  NAND2_X2 U1675 ( .A1(net155732), .A2(net155863), .ZN(net155782) );
  INV_X8 U1676 ( .A(net153819), .ZN(net155865) );
  NAND3_X2 U1677 ( .A1(net155493), .A2(net155865), .A3(net157351), .ZN(
        net155490) );
  NAND2_X2 U1678 ( .A1(net155496), .A2(net155865), .ZN(net155489) );
  NAND2_X4 U1679 ( .A1(y[2]), .A2(net155041), .ZN(net153819) );
  AOI21_X4 U1680 ( .B1(net153698), .B2(net157074), .A(net153700), .ZN(
        net153535) );
  NOR3_X4 U1681 ( .A1(net153960), .A2(net153961), .A3(net153962), .ZN(
        net153959) );
  OAI21_X4 U1682 ( .B1(n710), .B2(n782), .A(net153701), .ZN(net153699) );
  NAND2_X2 U1683 ( .A1(net153968), .A2(net153967), .ZN(n782) );
  NAND2_X4 U1684 ( .A1(n703), .A2(net153968), .ZN(net154356) );
  NAND3_X2 U1685 ( .A1(net154842), .A2(net154560), .A3(net153968), .ZN(
        net154773) );
  XNOR2_X2 U1686 ( .A(n696), .B(net156089), .ZN(net153952) );
  NAND2_X2 U1687 ( .A1(net154186), .A2(net154187), .ZN(net154171) );
  XNOR2_X2 U1688 ( .A(net154752), .B(net156169), .ZN(net157939) );
  NOR2_X4 U1689 ( .A1(net154744), .A2(net154745), .ZN(net154742) );
  INV_X4 U1690 ( .A(net154745), .ZN(net154701) );
  NAND4_X2 U1691 ( .A1(n2866), .A2(net153951), .A3(net153788), .A4(net153540), 
        .ZN(net154001) );
  NAND2_X1 U1692 ( .A1(net153547), .A2(net153951), .ZN(net154166) );
  NAND3_X2 U1693 ( .A1(net153951), .A2(net153780), .A3(net153540), .ZN(
        net153779) );
  NAND2_X4 U1694 ( .A1(net153952), .A2(net153953), .ZN(net153543) );
  INV_X8 U1695 ( .A(net157127), .ZN(net156089) );
  XNOR2_X2 U1696 ( .A(net154247), .B(n783), .ZN(net157127) );
  INV_X4 U1697 ( .A(n784), .ZN(n783) );
  XNOR2_X2 U1698 ( .A(n590), .B(n785), .ZN(n784) );
  INV_X4 U1699 ( .A(net154234), .ZN(n785) );
  OAI21_X4 U1700 ( .B1(net155885), .B2(net154852), .A(n786), .ZN(net154736) );
  NAND3_X2 U1701 ( .A1(net156073), .A2(net154795), .A3(net154796), .ZN(n786)
         );
  NOR3_X4 U1702 ( .A1(net153777), .A2(net153779), .A3(net153778), .ZN(
        net153673) );
  NOR2_X2 U1703 ( .A1(n589), .A2(net153977), .ZN(net153975) );
  NAND2_X2 U1704 ( .A1(net154323), .A2(net154322), .ZN(net154442) );
  NAND3_X2 U1705 ( .A1(n787), .A2(n788), .A3(n789), .ZN(net154328) );
  INV_X8 U1706 ( .A(net154477), .ZN(n791) );
  NAND3_X2 U1707 ( .A1(n791), .A2(net157527), .A3(net157773), .ZN(net154479)
         );
  NAND4_X1 U1708 ( .A1(n791), .A2(net153996), .A3(n792), .A4(net154341), .ZN(
        n787) );
  NAND2_X1 U1709 ( .A1(n791), .A2(net156869), .ZN(net154480) );
  NAND4_X1 U1710 ( .A1(net154332), .A2(net153996), .A3(n790), .A4(net154334), 
        .ZN(n789) );
  NOR3_X2 U1711 ( .A1(net154588), .A2(net154589), .A3(net156708), .ZN(n792) );
  INV_X2 U1712 ( .A(net153673), .ZN(net157619) );
  NAND2_X4 U1713 ( .A1(n796), .A2(n797), .ZN(n799) );
  INV_X1 U1714 ( .A(net153631), .ZN(n797) );
  INV_X4 U1715 ( .A(net153781), .ZN(n796) );
  NAND2_X1 U1716 ( .A1(net153631), .A2(net153781), .ZN(n798) );
  NAND2_X2 U1717 ( .A1(net158256), .A2(net153541), .ZN(net153777) );
  NAND2_X1 U1718 ( .A1(net153633), .A2(n794), .ZN(net153631) );
  XNOR2_X2 U1719 ( .A(net153630), .B(net153631), .ZN(net153517) );
  INV_X8 U1720 ( .A(n793), .ZN(n794) );
  XNOR2_X1 U1721 ( .A(n794), .B(n795), .ZN(net153743) );
  NAND2_X1 U1722 ( .A1(n794), .A2(n2809), .ZN(net156541) );
  NAND2_X4 U1723 ( .A1(net153856), .A2(n794), .ZN(net153863) );
  XNOR2_X2 U1724 ( .A(net156711), .B(net154006), .ZN(n793) );
  NOR2_X4 U1725 ( .A1(net153784), .A2(n795), .ZN(net153781) );
  INV_X4 U1726 ( .A(net153633), .ZN(n795) );
  XNOR2_X2 U1727 ( .A(net154531), .B(n800), .ZN(net154529) );
  NAND2_X2 U1728 ( .A1(net154533), .A2(net154534), .ZN(n800) );
  NAND2_X4 U1729 ( .A1(net154622), .A2(net154623), .ZN(net154537) );
  NAND2_X1 U1730 ( .A1(n2520), .A2(net156181), .ZN(net154687) );
  NAND2_X4 U1731 ( .A1(net154537), .A2(net154291), .ZN(net154033) );
  XNOR2_X2 U1732 ( .A(net156462), .B(net154786), .ZN(net154533) );
  INV_X4 U1733 ( .A(net154533), .ZN(net156664) );
  NAND2_X2 U1734 ( .A1(net156110), .A2(net154033), .ZN(net154151) );
  NAND2_X4 U1735 ( .A1(net157575), .A2(net157576), .ZN(net157578) );
  INV_X8 U1736 ( .A(net155820), .ZN(net155777) );
  AOI21_X2 U1737 ( .B1(n2042), .B2(n2066), .A(n2041), .ZN(n2045) );
  XNOR2_X2 U1738 ( .A(n1853), .B(n1852), .ZN(n801) );
  XNOR2_X2 U1739 ( .A(n807), .B(n1819), .ZN(n1852) );
  NOR2_X2 U1740 ( .A1(net153876), .A2(n2633), .ZN(n2636) );
  NAND2_X4 U1741 ( .A1(n2151), .A2(net156156), .ZN(n1073) );
  INV_X2 U1742 ( .A(net154687), .ZN(net154575) );
  INV_X4 U1743 ( .A(n2127), .ZN(n2147) );
  NOR2_X2 U1744 ( .A1(net154575), .A2(n2078), .ZN(n2079) );
  INV_X2 U1745 ( .A(n1772), .ZN(n802) );
  INV_X4 U1746 ( .A(n802), .ZN(n803) );
  OAI21_X1 U1747 ( .B1(n2896), .B2(n2895), .A(n2894), .ZN(n2901) );
  INV_X4 U1748 ( .A(n2217), .ZN(n1038) );
  NAND2_X2 U1749 ( .A1(n2217), .A2(n804), .ZN(n1040) );
  NAND2_X2 U1750 ( .A1(net154180), .A2(n2517), .ZN(net154320) );
  XNOR2_X2 U1751 ( .A(n2195), .B(n2194), .ZN(n804) );
  NOR3_X2 U1752 ( .A1(n606), .A2(n1167), .A3(net154061), .ZN(n2527) );
  INV_X1 U1753 ( .A(n1167), .ZN(n1064) );
  NAND2_X2 U1754 ( .A1(n1096), .A2(n1097), .ZN(n805) );
  NAND2_X4 U1755 ( .A1(net156663), .A2(net156664), .ZN(n1097) );
  INV_X1 U1756 ( .A(n1895), .ZN(n806) );
  INV_X4 U1757 ( .A(n1149), .ZN(n1577) );
  NAND2_X2 U1758 ( .A1(n1438), .A2(n1149), .ZN(n1667) );
  XNOR2_X2 U1759 ( .A(n2403), .B(n2402), .ZN(n809) );
  INV_X4 U1760 ( .A(net158330), .ZN(net154091) );
  XNOR2_X2 U1761 ( .A(n811), .B(n1256), .ZN(n810) );
  INV_X4 U1762 ( .A(n810), .ZN(n941) );
  XNOR2_X2 U1763 ( .A(n1255), .B(n1262), .ZN(n811) );
  INV_X4 U1764 ( .A(net153613), .ZN(net156130) );
  XNOR2_X2 U1765 ( .A(net156711), .B(net154006), .ZN(n812) );
  INV_X8 U1766 ( .A(net154667), .ZN(net156180) );
  NAND2_X4 U1767 ( .A1(n2609), .A2(n2611), .ZN(n2411) );
  INV_X2 U1768 ( .A(n1223), .ZN(n813) );
  NAND2_X2 U1769 ( .A1(n1655), .A2(n1657), .ZN(n1807) );
  INV_X2 U1770 ( .A(n1473), .ZN(n814) );
  INV_X4 U1771 ( .A(n1745), .ZN(n816) );
  NAND2_X4 U1772 ( .A1(n2138), .A2(n2142), .ZN(n2145) );
  NOR2_X4 U1773 ( .A1(n1857), .A2(n1858), .ZN(n817) );
  INV_X4 U1774 ( .A(n817), .ZN(n2027) );
  NAND2_X4 U1775 ( .A1(n2503), .A2(n2502), .ZN(n818) );
  NAND2_X4 U1776 ( .A1(n877), .A2(n878), .ZN(n2503) );
  NAND2_X4 U1777 ( .A1(n2453), .A2(n2452), .ZN(n2475) );
  OAI21_X2 U1778 ( .B1(n2451), .B2(n2483), .A(n2450), .ZN(n2452) );
  NOR2_X4 U1779 ( .A1(x[2]), .A2(x[1]), .ZN(n1444) );
  BUF_X8 U1780 ( .A(n572), .Z(n821) );
  XOR2_X1 U1781 ( .A(n1043), .B(n1914), .Z(n822) );
  NAND2_X2 U1782 ( .A1(n2385), .A2(n2499), .ZN(n2430) );
  NAND2_X4 U1783 ( .A1(n1200), .A2(n1199), .ZN(n1287) );
  NAND2_X2 U1784 ( .A1(n915), .A2(n2514), .ZN(n1761) );
  INV_X8 U1785 ( .A(n1897), .ZN(n1996) );
  INV_X4 U1786 ( .A(n2808), .ZN(n2654) );
  NOR2_X2 U1787 ( .A1(n1136), .A2(n1137), .ZN(n1138) );
  XNOR2_X2 U1788 ( .A(n1843), .B(n1842), .ZN(n824) );
  INV_X8 U1789 ( .A(n2631), .ZN(net158270) );
  NAND2_X4 U1790 ( .A1(n2626), .A2(n2625), .ZN(net158266) );
  INV_X8 U1791 ( .A(n2624), .ZN(n2626) );
  INV_X8 U1792 ( .A(n1814), .ZN(n1751) );
  XNOR2_X1 U1793 ( .A(n2543), .B(net153743), .ZN(n2728) );
  INV_X8 U1794 ( .A(net156130), .ZN(net157527) );
  NAND2_X4 U1795 ( .A1(n2582), .A2(n2581), .ZN(net158256) );
  NAND3_X1 U1796 ( .A1(n2505), .A2(net153835), .A3(net153829), .ZN(n2486) );
  NOR2_X2 U1797 ( .A1(net154169), .A2(net153550), .ZN(n2420) );
  XNOR2_X1 U1798 ( .A(n1879), .B(net155057), .ZN(n1816) );
  OAI22_X1 U1799 ( .A1(n2705), .A2(net154784), .B1(net155835), .B2(n2013), 
        .ZN(n2022) );
  NAND2_X1 U1800 ( .A1(n841), .A2(net156180), .ZN(n838) );
  NAND2_X4 U1801 ( .A1(n2509), .A2(n2658), .ZN(n2510) );
  NOR2_X2 U1802 ( .A1(n2110), .A2(n2178), .ZN(n2062) );
  NOR2_X2 U1803 ( .A1(net156130), .A2(n805), .ZN(n826) );
  INV_X1 U1804 ( .A(net153937), .ZN(net158242) );
  INV_X8 U1805 ( .A(n1856), .ZN(n1857) );
  INV_X1 U1806 ( .A(net157381), .ZN(net154971) );
  XNOR2_X1 U1807 ( .A(n2786), .B(n2653), .ZN(n828) );
  NAND4_X2 U1808 ( .A1(n2408), .A2(n2409), .A3(n2456), .A4(n2370), .ZN(n2410)
         );
  INV_X8 U1809 ( .A(n2206), .ZN(n1021) );
  XNOR2_X2 U1810 ( .A(n1914), .B(n1931), .ZN(n830) );
  NAND2_X4 U1811 ( .A1(n1027), .A2(n570), .ZN(n863) );
  NAND2_X4 U1812 ( .A1(x[13]), .A2(n2606), .ZN(n1705) );
  NAND2_X2 U1813 ( .A1(n2824), .A2(n2644), .ZN(n2692) );
  NAND2_X2 U1814 ( .A1(n2273), .A2(n944), .ZN(n2308) );
  INV_X2 U1815 ( .A(n1889), .ZN(n831) );
  BUF_X32 U1816 ( .A(n1430), .Z(n832) );
  XNOR2_X2 U1817 ( .A(n886), .B(n1021), .ZN(n833) );
  INV_X1 U1818 ( .A(n1501), .ZN(n834) );
  INV_X8 U1819 ( .A(n1833), .ZN(n1804) );
  XNOR2_X2 U1820 ( .A(n1241), .B(x[5]), .ZN(n836) );
  XNOR2_X2 U1821 ( .A(n2554), .B(n2560), .ZN(net153977) );
  NAND2_X2 U1822 ( .A1(n806), .A2(n825), .ZN(n1872) );
  NAND2_X2 U1823 ( .A1(n1125), .A2(n1992), .ZN(n1995) );
  INV_X2 U1824 ( .A(n1888), .ZN(n837) );
  NAND2_X2 U1825 ( .A1(n2050), .A2(net158130), .ZN(net154734) );
  NAND2_X4 U1826 ( .A1(n1905), .A2(n1971), .ZN(net154877) );
  INV_X8 U1827 ( .A(n1580), .ZN(n839) );
  INV_X4 U1828 ( .A(n2154), .ZN(n840) );
  INV_X8 U1829 ( .A(net154025), .ZN(n841) );
  INV_X8 U1830 ( .A(net154956), .ZN(net156405) );
  INV_X2 U1831 ( .A(n1573), .ZN(n842) );
  INV_X1 U1832 ( .A(n543), .ZN(n843) );
  INV_X2 U1833 ( .A(n2232), .ZN(n2372) );
  INV_X2 U1834 ( .A(n1370), .ZN(n844) );
  INV_X4 U1835 ( .A(n1935), .ZN(n1043) );
  OAI22_X4 U1836 ( .A1(n1175), .A2(n2469), .B1(n2686), .B2(net155869), .ZN(
        n846) );
  OAI21_X1 U1837 ( .B1(n829), .B2(net155869), .A(n1568), .ZN(n847) );
  XNOR2_X1 U1838 ( .A(n1236), .B(n1235), .ZN(n848) );
  INV_X4 U1839 ( .A(net156708), .ZN(net158146) );
  NAND2_X1 U1840 ( .A1(n836), .A2(n542), .ZN(n1291) );
  XNOR2_X2 U1841 ( .A(n1241), .B(x[5]), .ZN(n849) );
  CLKBUF_X3 U1842 ( .A(n2678), .Z(n850) );
  INV_X8 U1843 ( .A(n2891), .ZN(n852) );
  INV_X8 U1844 ( .A(n2890), .ZN(n2891) );
  INV_X2 U1845 ( .A(n1099), .ZN(n1145) );
  NAND2_X4 U1846 ( .A1(n1398), .A2(n1397), .ZN(n1376) );
  NAND2_X4 U1847 ( .A1(n2877), .A2(n2876), .ZN(net158121) );
  INV_X4 U1848 ( .A(net158116), .ZN(net158117) );
  NAND2_X2 U1849 ( .A1(n2918), .A2(n2917), .ZN(n1121) );
  NAND2_X4 U1850 ( .A1(n1618), .A2(n1684), .ZN(n1593) );
  XNOR2_X1 U1851 ( .A(n629), .B(n1232), .ZN(n1237) );
  XNOR2_X2 U1852 ( .A(n2726), .B(n2727), .ZN(n854) );
  NAND2_X4 U1853 ( .A1(n2724), .A2(n2725), .ZN(n2726) );
  NAND2_X2 U1854 ( .A1(n841), .A2(n2522), .ZN(n2523) );
  INV_X8 U1855 ( .A(n856), .ZN(n857) );
  INV_X4 U1856 ( .A(n2535), .ZN(n1053) );
  OAI21_X1 U1857 ( .B1(n1495), .B2(n564), .A(n539), .ZN(n1499) );
  NOR2_X2 U1858 ( .A1(n1783), .A2(n1442), .ZN(net155493) );
  AOI21_X2 U1859 ( .B1(n1961), .B2(n580), .A(net154760), .ZN(n1962) );
  NOR2_X2 U1860 ( .A1(n1963), .A2(n1962), .ZN(n1984) );
  NAND2_X2 U1861 ( .A1(n2565), .A2(net153545), .ZN(net153962) );
  NAND2_X1 U1862 ( .A1(net154025), .A2(n2065), .ZN(n2018) );
  NAND2_X2 U1863 ( .A1(n2065), .A2(net154025), .ZN(n2002) );
  AOI21_X2 U1864 ( .B1(n2252), .B2(n2253), .A(n2251), .ZN(n2254) );
  NAND2_X4 U1865 ( .A1(n2606), .A2(n516), .ZN(n1382) );
  INV_X4 U1866 ( .A(n899), .ZN(n858) );
  AND2_X4 U1867 ( .A1(n2316), .A2(n2552), .ZN(n859) );
  NAND3_X1 U1868 ( .A1(n2325), .A2(net154349), .A3(n2324), .ZN(n2872) );
  INV_X1 U1869 ( .A(n1009), .ZN(n947) );
  XOR2_X2 U1870 ( .A(n2618), .B(n565), .Z(n860) );
  OAI22_X2 U1871 ( .A1(net155885), .A2(n2469), .B1(net155857), .B2(n545), .ZN(
        n2618) );
  XNOR2_X1 U1872 ( .A(n2562), .B(net153975), .ZN(n861) );
  INV_X2 U1873 ( .A(net154250), .ZN(net158084) );
  NAND2_X4 U1874 ( .A1(n1837), .A2(n1836), .ZN(net157381) );
  XNOR2_X2 U1875 ( .A(n1484), .B(x[11]), .ZN(n862) );
  INV_X4 U1876 ( .A(n2004), .ZN(n2008) );
  NAND2_X4 U1877 ( .A1(n2017), .A2(n2002), .ZN(n2269) );
  NAND2_X2 U1878 ( .A1(n1213), .A2(n1116), .ZN(n1239) );
  NAND2_X2 U1879 ( .A1(n1060), .A2(n2851), .ZN(n2791) );
  INV_X2 U1880 ( .A(n1016), .ZN(n2226) );
  INV_X4 U1881 ( .A(n1994), .ZN(n1850) );
  NAND2_X4 U1882 ( .A1(n817), .A2(n1859), .ZN(n1862) );
  NOR2_X2 U1883 ( .A1(n1735), .A2(n1734), .ZN(n1739) );
  OAI221_X2 U1884 ( .B1(n2631), .B2(net153829), .C1(n2631), .C2(n679), .A(
        n2630), .ZN(n2632) );
  NAND2_X2 U1885 ( .A1(n1280), .A2(n864), .ZN(n866) );
  INV_X2 U1886 ( .A(n1283), .ZN(n864) );
  NAND2_X2 U1887 ( .A1(n1254), .A2(n1253), .ZN(n869) );
  NAND2_X4 U1888 ( .A1(n867), .A2(n868), .ZN(n870) );
  NAND2_X4 U1889 ( .A1(n869), .A2(n870), .ZN(n1343) );
  INV_X4 U1890 ( .A(n1254), .ZN(n867) );
  INV_X4 U1891 ( .A(n1253), .ZN(n868) );
  NAND2_X4 U1892 ( .A1(n1243), .A2(n1242), .ZN(n1283) );
  NAND2_X2 U1893 ( .A1(n1252), .A2(n1251), .ZN(n1253) );
  NAND2_X2 U1894 ( .A1(n1690), .A2(n1689), .ZN(n873) );
  NAND2_X4 U1895 ( .A1(n871), .A2(n872), .ZN(n874) );
  NAND2_X4 U1896 ( .A1(n873), .A2(n874), .ZN(n1733) );
  INV_X4 U1897 ( .A(n1690), .ZN(n871) );
  INV_X4 U1898 ( .A(n1689), .ZN(n872) );
  INV_X2 U1899 ( .A(n1733), .ZN(n1734) );
  NAND2_X2 U1900 ( .A1(n875), .A2(n876), .ZN(n878) );
  INV_X1 U1901 ( .A(n2616), .ZN(n876) );
  INV_X2 U1902 ( .A(net153856), .ZN(net153853) );
  INV_X4 U1903 ( .A(n2642), .ZN(n2628) );
  NAND2_X4 U1904 ( .A1(n879), .A2(n880), .ZN(n882) );
  INV_X4 U1905 ( .A(n2315), .ZN(n879) );
  INV_X16 U1906 ( .A(net153818), .ZN(net155884) );
  INV_X8 U1907 ( .A(net154885), .ZN(net154308) );
  INV_X1 U1908 ( .A(n2329), .ZN(n2078) );
  NAND2_X1 U1909 ( .A1(n2096), .A2(n2329), .ZN(n2102) );
  NOR2_X4 U1910 ( .A1(n1175), .A2(net154940), .ZN(n1924) );
  INV_X8 U1911 ( .A(n2550), .ZN(n883) );
  NAND2_X4 U1912 ( .A1(n1206), .A2(n1205), .ZN(n1232) );
  INV_X4 U1913 ( .A(n1232), .ZN(n1234) );
  AOI21_X2 U1914 ( .B1(n1575), .B2(n1574), .A(n1573), .ZN(n1576) );
  CLKBUF_X3 U1915 ( .A(net154699), .Z(net157644) );
  OAI21_X2 U1916 ( .B1(n803), .B2(n915), .A(n1061), .ZN(n1766) );
  XNOR2_X2 U1917 ( .A(n1853), .B(n1852), .ZN(n2028) );
  NAND2_X4 U1918 ( .A1(n1583), .A2(n932), .ZN(n1578) );
  OR2_X2 U1919 ( .A1(n2547), .A2(n2548), .ZN(n1085) );
  XNOR2_X2 U1920 ( .A(net154031), .B(n2277), .ZN(n2271) );
  NAND2_X4 U1921 ( .A1(n884), .A2(x[14]), .ZN(n885) );
  NAND2_X4 U1922 ( .A1(n1716), .A2(n885), .ZN(n1746) );
  INV_X1 U1923 ( .A(n1174), .ZN(n884) );
  NAND2_X2 U1924 ( .A1(n928), .A2(n929), .ZN(n2696) );
  NOR3_X2 U1925 ( .A1(n1739), .A2(n1738), .A3(n1737), .ZN(n1742) );
  NAND2_X1 U1926 ( .A1(net153784), .A2(n812), .ZN(n928) );
  NAND2_X4 U1927 ( .A1(n1200), .A2(n1199), .ZN(n1186) );
  NAND2_X4 U1928 ( .A1(n2390), .A2(n2389), .ZN(n886) );
  INV_X2 U1929 ( .A(n2077), .ZN(n2000) );
  NAND2_X4 U1930 ( .A1(n1972), .A2(n1973), .ZN(n1845) );
  NAND2_X4 U1931 ( .A1(n2081), .A2(n805), .ZN(n2097) );
  NOR4_X4 U1932 ( .A1(x[6]), .A2(x[5]), .A3(x[8]), .A4(x[7]), .ZN(n887) );
  NAND2_X2 U1933 ( .A1(n606), .A2(n2435), .ZN(n890) );
  NAND2_X4 U1934 ( .A1(n888), .A2(n889), .ZN(n891) );
  INV_X4 U1935 ( .A(n2435), .ZN(n888) );
  INV_X4 U1936 ( .A(net153835), .ZN(net153833) );
  OAI21_X4 U1937 ( .B1(n2300), .B2(n2299), .A(n2298), .ZN(n2310) );
  INV_X4 U1938 ( .A(n2575), .ZN(n2357) );
  NAND2_X2 U1939 ( .A1(n1610), .A2(n546), .ZN(n892) );
  NAND2_X4 U1940 ( .A1(n892), .A2(n893), .ZN(n1147) );
  XNOR2_X2 U1941 ( .A(n872), .B(n1735), .ZN(n1611) );
  NAND2_X2 U1942 ( .A1(n894), .A2(n895), .ZN(n896) );
  NAND2_X4 U1943 ( .A1(n896), .A2(n2220), .ZN(n2224) );
  INV_X2 U1944 ( .A(n2218), .ZN(n894) );
  NAND2_X4 U1945 ( .A1(n1160), .A2(n1159), .ZN(n2562) );
  NOR2_X4 U1946 ( .A1(x[7]), .A2(x[8]), .ZN(net157892) );
  INV_X4 U1947 ( .A(n1878), .ZN(n897) );
  INV_X4 U1948 ( .A(n1878), .ZN(n1883) );
  BUF_X8 U1949 ( .A(n1795), .Z(n899) );
  INV_X1 U1950 ( .A(n1881), .ZN(n1774) );
  NOR2_X4 U1951 ( .A1(n2883), .A2(n2882), .ZN(n2884) );
  NOR2_X4 U1952 ( .A1(n1469), .A2(n1468), .ZN(n1478) );
  INV_X8 U1953 ( .A(n1657), .ZN(n1580) );
  NAND2_X4 U1954 ( .A1(n1528), .A2(n1527), .ZN(n1530) );
  NAND3_X2 U1955 ( .A1(n2716), .A2(n2909), .A3(n2715), .ZN(n2894) );
  INV_X8 U1956 ( .A(n1886), .ZN(n1795) );
  NAND2_X2 U1957 ( .A1(n1380), .A2(n1338), .ZN(n903) );
  NAND2_X4 U1958 ( .A1(n901), .A2(n902), .ZN(n904) );
  NAND2_X4 U1959 ( .A1(n903), .A2(n904), .ZN(n1365) );
  INV_X2 U1960 ( .A(n1380), .ZN(n901) );
  INV_X4 U1961 ( .A(n1338), .ZN(n902) );
  NAND2_X2 U1962 ( .A1(n1282), .A2(x[5]), .ZN(n906) );
  NAND2_X4 U1963 ( .A1(n905), .A2(net157848), .ZN(n907) );
  NAND2_X4 U1964 ( .A1(n907), .A2(n906), .ZN(n1148) );
  INV_X4 U1965 ( .A(n1282), .ZN(n905) );
  INV_X4 U1966 ( .A(x[5]), .ZN(net157848) );
  NAND2_X4 U1967 ( .A1(n1621), .A2(n1620), .ZN(n1638) );
  NAND2_X2 U1968 ( .A1(net154620), .A2(net154621), .ZN(net157577) );
  INV_X1 U1969 ( .A(n1320), .ZN(n1278) );
  NAND2_X2 U1970 ( .A1(n1034), .A2(n1033), .ZN(n1036) );
  NAND2_X2 U1971 ( .A1(net155315), .A2(n1787), .ZN(n1779) );
  NOR2_X2 U1972 ( .A1(n2379), .A2(n2368), .ZN(n2369) );
  INV_X2 U1973 ( .A(n2720), .ZN(n1028) );
  NAND2_X1 U1974 ( .A1(n1546), .A2(n843), .ZN(n1613) );
  INV_X4 U1975 ( .A(n2518), .ZN(n908) );
  INV_X4 U1976 ( .A(n2665), .ZN(n2518) );
  INV_X4 U1977 ( .A(n2352), .ZN(n2356) );
  NAND4_X4 U1978 ( .A1(net154943), .A2(net155315), .A3(n1417), .A4(net157892), 
        .ZN(n1418) );
  NAND2_X4 U1979 ( .A1(n1572), .A2(net155873), .ZN(n1574) );
  NOR3_X4 U1980 ( .A1(n1672), .A2(n1673), .A3(n1671), .ZN(n909) );
  NAND2_X2 U1981 ( .A1(n1669), .A2(n1668), .ZN(n911) );
  INV_X1 U1982 ( .A(n1665), .ZN(n1669) );
  XNOR2_X2 U1983 ( .A(n1902), .B(net154968), .ZN(n1846) );
  INV_X4 U1984 ( .A(n1127), .ZN(n975) );
  NAND3_X2 U1985 ( .A1(n2894), .A2(n2898), .A3(n2890), .ZN(n2850) );
  NAND2_X4 U1986 ( .A1(n1247), .A2(n1256), .ZN(n1406) );
  NAND2_X4 U1987 ( .A1(net157767), .A2(net156110), .ZN(n913) );
  NAND2_X4 U1988 ( .A1(net157769), .A2(n913), .ZN(n944) );
  INV_X4 U1989 ( .A(net154660), .ZN(net157767) );
  INV_X4 U1990 ( .A(n1826), .ZN(n1874) );
  NAND2_X4 U1991 ( .A1(n2438), .A2(n2584), .ZN(n2496) );
  NAND2_X1 U1992 ( .A1(n2174), .A2(n2308), .ZN(n2105) );
  NAND2_X4 U1993 ( .A1(n1479), .A2(n1546), .ZN(n1480) );
  INV_X8 U1994 ( .A(n948), .ZN(n949) );
  NAND2_X4 U1995 ( .A1(n1446), .A2(n1445), .ZN(n948) );
  NOR2_X4 U1996 ( .A1(x[8]), .A2(x[7]), .ZN(n1445) );
  NAND2_X2 U1997 ( .A1(net153835), .A2(net153829), .ZN(n2507) );
  INV_X1 U1998 ( .A(n2308), .ZN(n2179) );
  NAND2_X1 U1999 ( .A1(n2103), .A2(n2308), .ZN(n2104) );
  INV_X2 U2000 ( .A(n2175), .ZN(n2165) );
  NOR2_X4 U2001 ( .A1(n2639), .A2(n2638), .ZN(n2640) );
  INV_X4 U2002 ( .A(n1442), .ZN(n914) );
  CLKBUF_X2 U2003 ( .A(n2337), .Z(n915) );
  INV_X4 U2004 ( .A(n1264), .ZN(n1267) );
  NAND2_X4 U2005 ( .A1(n501), .A2(n1864), .ZN(n1854) );
  NOR2_X2 U2006 ( .A1(n2232), .A2(n917), .ZN(n916) );
  OAI21_X4 U2007 ( .B1(n1384), .B2(n1383), .A(n823), .ZN(n1393) );
  NAND2_X2 U2008 ( .A1(n517), .A2(n1907), .ZN(n1908) );
  NAND2_X4 U2009 ( .A1(n1826), .A2(n1828), .ZN(n1853) );
  NOR2_X2 U2010 ( .A1(n898), .A2(n1772), .ZN(n1773) );
  NAND2_X2 U2011 ( .A1(n1611), .A2(n1612), .ZN(n986) );
  NAND3_X4 U2012 ( .A1(n1841), .A2(n1904), .A3(n1916), .ZN(n1843) );
  NAND3_X2 U2013 ( .A1(n2369), .A2(n2370), .A3(n2454), .ZN(n2374) );
  NOR2_X2 U2014 ( .A1(n2288), .A2(n2172), .ZN(n2036) );
  NAND2_X2 U2015 ( .A1(n535), .A2(n1780), .ZN(n1786) );
  NOR2_X2 U2016 ( .A1(x[4]), .A2(x[15]), .ZN(n1782) );
  INV_X2 U2017 ( .A(n1028), .ZN(n1029) );
  NAND2_X1 U2018 ( .A1(n570), .A2(n1027), .ZN(net154589) );
  INV_X2 U2019 ( .A(net153796), .ZN(net153671) );
  OAI21_X4 U2020 ( .B1(x[9]), .B2(net156405), .A(x[10]), .ZN(n1546) );
  NOR2_X2 U2021 ( .A1(net154575), .A2(n2155), .ZN(n2156) );
  NAND2_X2 U2022 ( .A1(n2082), .A2(net154687), .ZN(n2301) );
  OAI21_X2 U2023 ( .B1(n1467), .B2(net155869), .A(n1466), .ZN(n1655) );
  NAND2_X1 U2024 ( .A1(n1459), .A2(n633), .ZN(n1630) );
  NAND2_X2 U2025 ( .A1(n1827), .A2(n1816), .ZN(n1128) );
  AND2_X2 U2026 ( .A1(n1410), .A2(n1404), .ZN(n921) );
  NAND2_X4 U2027 ( .A1(n2554), .A2(n2553), .ZN(n1163) );
  INV_X8 U2028 ( .A(n2533), .ZN(n1172) );
  INV_X1 U2029 ( .A(n2697), .ZN(n2437) );
  NAND2_X2 U2030 ( .A1(n1275), .A2(n1273), .ZN(n924) );
  NAND2_X2 U2031 ( .A1(n922), .A2(n923), .ZN(n925) );
  INV_X4 U2032 ( .A(n1275), .ZN(n922) );
  NAND2_X4 U2033 ( .A1(x[1]), .A2(x[0]), .ZN(n926) );
  NAND2_X4 U2034 ( .A1(net157664), .A2(net157665), .ZN(n927) );
  NAND2_X4 U2035 ( .A1(n926), .A2(n927), .ZN(net155787) );
  INV_X8 U2036 ( .A(x[1]), .ZN(net157664) );
  INV_X32 U2037 ( .A(x[0]), .ZN(net157665) );
  OAI21_X4 U2038 ( .B1(net155787), .B2(n1559), .A(net155799), .ZN(n1286) );
  INV_X4 U2039 ( .A(n2703), .ZN(n1034) );
  XNOR2_X1 U2040 ( .A(n832), .B(n602), .ZN(n1428) );
  NAND2_X2 U2041 ( .A1(net157651), .A2(n2767), .ZN(n929) );
  INV_X2 U2042 ( .A(net153784), .ZN(net157651) );
  INV_X2 U2043 ( .A(n1969), .ZN(n1010) );
  INV_X4 U2044 ( .A(net154621), .ZN(net157576) );
  OAI21_X1 U2045 ( .B1(net155827), .B2(n1763), .A(n1762), .ZN(n1855) );
  OAI22_X1 U2046 ( .A1(net155896), .A2(net155324), .B1(net155841), .B2(n1763), 
        .ZN(n1728) );
  NAND2_X4 U2047 ( .A1(n2113), .A2(n2205), .ZN(n2116) );
  INV_X2 U2048 ( .A(net156089), .ZN(net154083) );
  NAND2_X2 U2049 ( .A1(n1150), .A2(n1576), .ZN(n982) );
  NAND2_X4 U2050 ( .A1(net153541), .A2(net158256), .ZN(n2698) );
  INV_X4 U2051 ( .A(n1667), .ZN(n931) );
  INV_X8 U2052 ( .A(n931), .ZN(n932) );
  INV_X2 U2053 ( .A(n933), .ZN(n934) );
  NOR2_X4 U2054 ( .A1(n1413), .A2(net155869), .ZN(n1373) );
  NAND2_X2 U2055 ( .A1(net157619), .A2(n935), .ZN(n936) );
  NAND2_X2 U2056 ( .A1(n936), .A2(n677), .ZN(n2700) );
  NAND3_X2 U2057 ( .A1(y[0]), .A2(net155041), .A3(x[3]), .ZN(n1214) );
  NOR2_X4 U2058 ( .A1(x[4]), .A2(x[3]), .ZN(n1446) );
  NAND2_X4 U2059 ( .A1(net155513), .A2(net155514), .ZN(net157615) );
  INV_X32 U2060 ( .A(x[6]), .ZN(net155514) );
  NAND2_X4 U2061 ( .A1(n938), .A2(n601), .ZN(net154158) );
  NAND2_X4 U2062 ( .A1(n1887), .A2(n858), .ZN(n1890) );
  OAI21_X2 U2063 ( .B1(n1888), .B2(n899), .A(n1752), .ZN(n1753) );
  INV_X1 U2064 ( .A(n1220), .ZN(n1193) );
  INV_X4 U2065 ( .A(n1567), .ZN(n1723) );
  NOR2_X4 U2066 ( .A1(n918), .A2(n1482), .ZN(n1484) );
  INV_X1 U2067 ( .A(n1767), .ZN(n1681) );
  INV_X4 U2068 ( .A(n1569), .ZN(n1131) );
  XNOR2_X2 U2069 ( .A(n940), .B(n1593), .ZN(n939) );
  NAND3_X2 U2070 ( .A1(net155315), .A2(n731), .A3(n1443), .ZN(n1840) );
  NAND2_X4 U2071 ( .A1(n1381), .A2(net155859), .ZN(n1397) );
  INV_X4 U2072 ( .A(net154356), .ZN(net154423) );
  INV_X4 U2073 ( .A(n1796), .ZN(n942) );
  INV_X4 U2074 ( .A(n1796), .ZN(n1831) );
  NOR2_X1 U2075 ( .A1(n2730), .A2(n2729), .ZN(n2735) );
  INV_X8 U2076 ( .A(net157404), .ZN(n943) );
  OAI22_X4 U2077 ( .A1(n1174), .A2(net154852), .B1(net155869), .B2(n2093), 
        .ZN(net154817) );
  NAND2_X2 U2078 ( .A1(n716), .A2(n718), .ZN(n2053) );
  OAI22_X4 U2079 ( .A1(net155885), .A2(n2057), .B1(n2212), .B2(net155857), 
        .ZN(n2115) );
  NAND2_X4 U2080 ( .A1(n2230), .A2(n2358), .ZN(n2472) );
  NAND2_X2 U2081 ( .A1(n2622), .A2(n819), .ZN(net156711) );
  INV_X2 U2082 ( .A(n2780), .ZN(n2751) );
  INV_X8 U2083 ( .A(n1746), .ZN(n1794) );
  INV_X4 U2084 ( .A(net157531), .ZN(net157532) );
  NOR2_X2 U2085 ( .A1(n1117), .A2(n1840), .ZN(n1841) );
  XNOR2_X2 U2086 ( .A(n1365), .B(n946), .ZN(n945) );
  INV_X4 U2087 ( .A(net154829), .ZN(net157542) );
  INV_X8 U2088 ( .A(net154682), .ZN(net154829) );
  INV_X4 U2089 ( .A(n1970), .ZN(n1009) );
  NOR2_X1 U2090 ( .A1(n1314), .A2(n532), .ZN(n1277) );
  INV_X8 U2091 ( .A(n2492), .ZN(n1063) );
  NAND3_X2 U2092 ( .A1(n1711), .A2(n1710), .A3(n1781), .ZN(n1712) );
  XNOR2_X2 U2093 ( .A(n1526), .B(n564), .ZN(n1528) );
  INV_X8 U2094 ( .A(n1791), .ZN(n1916) );
  INV_X16 U2095 ( .A(x[6]), .ZN(net157521) );
  INV_X4 U2096 ( .A(n1687), .ZN(n1005) );
  INV_X32 U2097 ( .A(x[4]), .ZN(net155665) );
  INV_X32 U2098 ( .A(x[4]), .ZN(net155645) );
  AOI21_X2 U2099 ( .B1(n1309), .B2(n1308), .A(n1307), .ZN(n1311) );
  INV_X8 U2100 ( .A(n2811), .ZN(n2722) );
  AOI21_X4 U2101 ( .B1(n1571), .B2(n932), .A(n1570), .ZN(n1579) );
  NOR2_X4 U2102 ( .A1(n2616), .A2(n809), .ZN(n2612) );
  INV_X2 U2103 ( .A(n2797), .ZN(n2799) );
  AOI21_X2 U2104 ( .B1(n2877), .B2(n2876), .A(n2875), .ZN(n2885) );
  INV_X8 U2105 ( .A(n1152), .ZN(n2207) );
  INV_X4 U2106 ( .A(net155314), .ZN(net155506) );
  NAND2_X4 U2107 ( .A1(n2614), .A2(n1055), .ZN(n2616) );
  NAND2_X4 U2108 ( .A1(n1053), .A2(n1054), .ZN(n1055) );
  XNOR2_X1 U2109 ( .A(n1950), .B(n1949), .ZN(n2290) );
  NAND2_X1 U2110 ( .A1(n841), .A2(n2080), .ZN(n950) );
  NAND3_X1 U2111 ( .A1(n2079), .A2(n951), .A3(n2187), .ZN(n2302) );
  INV_X4 U2112 ( .A(n950), .ZN(n951) );
  INV_X2 U2113 ( .A(n1797), .ZN(n1800) );
  NAND2_X4 U2114 ( .A1(n2054), .A2(net154728), .ZN(n2122) );
  NAND2_X1 U2115 ( .A1(n506), .A2(n2697), .ZN(n2422) );
  NOR2_X1 U2116 ( .A1(n2698), .A2(n2697), .ZN(n2495) );
  NAND2_X2 U2117 ( .A1(n2745), .A2(n2744), .ZN(n954) );
  INV_X4 U2118 ( .A(n2745), .ZN(n952) );
  INV_X1 U2119 ( .A(n2744), .ZN(n953) );
  NAND2_X4 U2120 ( .A1(n1880), .A2(n1879), .ZN(n1882) );
  NAND3_X4 U2121 ( .A1(net155775), .A2(net155773), .A3(net157440), .ZN(n956)
         );
  NAND2_X4 U2122 ( .A1(n2763), .A2(n2830), .ZN(n2842) );
  AOI21_X4 U2123 ( .B1(n1890), .B2(n1889), .A(n1888), .ZN(n1894) );
  NAND2_X4 U2124 ( .A1(n2350), .A2(n2515), .ZN(net153623) );
  NAND2_X2 U2125 ( .A1(n2492), .A2(n1167), .ZN(n1065) );
  NAND2_X4 U2126 ( .A1(n2350), .A2(n601), .ZN(n2478) );
  NAND2_X4 U2127 ( .A1(n581), .A2(n2571), .ZN(n2866) );
  INV_X4 U2128 ( .A(n2632), .ZN(n2637) );
  XNOR2_X2 U2129 ( .A(x[15]), .B(n1776), .ZN(n958) );
  NOR2_X2 U2130 ( .A1(n1899), .A2(n1898), .ZN(n1900) );
  NAND2_X4 U2131 ( .A1(n2739), .A2(n2770), .ZN(n2892) );
  NAND2_X4 U2132 ( .A1(n1504), .A2(n960), .ZN(n1539) );
  INV_X4 U2133 ( .A(n959), .ZN(n960) );
  INV_X32 U2134 ( .A(x[2]), .ZN(net157450) );
  INV_X32 U2135 ( .A(x[2]), .ZN(net157451) );
  XNOR2_X2 U2136 ( .A(n886), .B(n961), .ZN(net154339) );
  XOR2_X1 U2137 ( .A(n2206), .B(n2658), .Z(n961) );
  NAND2_X2 U2138 ( .A1(n1299), .A2(n1370), .ZN(n1301) );
  INV_X4 U2139 ( .A(n1651), .ZN(n1731) );
  NAND2_X4 U2140 ( .A1(n964), .A2(n965), .ZN(n2568) );
  INV_X2 U2141 ( .A(n2160), .ZN(n963) );
  NAND2_X1 U2142 ( .A1(n2303), .A2(n2159), .ZN(n2160) );
  INV_X32 U2143 ( .A(x[0]), .ZN(net157440) );
  OAI21_X4 U2144 ( .B1(n546), .B2(n712), .A(n851), .ZN(n1833) );
  XNOR2_X1 U2145 ( .A(n2062), .B(net158242), .ZN(result[22]) );
  NAND2_X2 U2146 ( .A1(n2045), .A2(n2044), .ZN(n2061) );
  OAI21_X2 U2147 ( .B1(n2070), .B2(n2020), .A(n2019), .ZN(n2021) );
  INV_X8 U2148 ( .A(n1462), .ZN(n1473) );
  NAND4_X2 U2149 ( .A1(n2867), .A2(n551), .A3(n686), .A4(net153543), .ZN(n2868) );
  INV_X8 U2150 ( .A(n2358), .ZN(n2359) );
  NOR2_X4 U2151 ( .A1(n1148), .A2(net155855), .ZN(n1329) );
  NAND2_X4 U2152 ( .A1(n966), .A2(n967), .ZN(net157424) );
  INV_X4 U2153 ( .A(net157424), .ZN(net154862) );
  INV_X32 U2154 ( .A(x[14]), .ZN(n966) );
  INV_X32 U2155 ( .A(x[13]), .ZN(n967) );
  NOR2_X4 U2156 ( .A1(n1379), .A2(n1378), .ZN(n1384) );
  NOR2_X2 U2157 ( .A1(n2732), .A2(n1022), .ZN(n2591) );
  INV_X2 U2158 ( .A(n2689), .ZN(n2732) );
  XNOR2_X2 U2159 ( .A(n1224), .B(n1290), .ZN(n1228) );
  OAI21_X4 U2160 ( .B1(n2494), .B2(n2493), .A(n2866), .ZN(n2438) );
  INV_X1 U2161 ( .A(net155508), .ZN(net157416) );
  INV_X32 U2162 ( .A(x[0]), .ZN(net155508) );
  NAND2_X2 U2163 ( .A1(n852), .A2(n2792), .ZN(n2794) );
  NAND2_X2 U2164 ( .A1(n2086), .A2(n2087), .ZN(n993) );
  INV_X4 U2165 ( .A(n2828), .ZN(n2893) );
  INV_X4 U2166 ( .A(n1941), .ZN(n1926) );
  OAI21_X2 U2167 ( .B1(net155839), .B2(n1937), .A(n1930), .ZN(n2335) );
  NOR4_X2 U2168 ( .A1(net155457), .A2(n649), .A3(n1598), .A4(n1597), .ZN(n1558) );
  INV_X4 U2169 ( .A(n2151), .ZN(n1072) );
  OAI211_X4 U2170 ( .C1(n2066), .C2(net158146), .A(n2523), .B(net157527), .ZN(
        n2815) );
  NAND2_X2 U2171 ( .A1(n2247), .A2(net154250), .ZN(n2381) );
  INV_X8 U2172 ( .A(n1827), .ZN(n1127) );
  INV_X8 U2173 ( .A(n1423), .ZN(n1441) );
  XNOR2_X2 U2174 ( .A(n1497), .B(n1496), .ZN(n1498) );
  NAND2_X4 U2175 ( .A1(net155696), .A2(net155665), .ZN(n968) );
  NAND2_X4 U2176 ( .A1(n1279), .A2(n1292), .ZN(n1244) );
  NAND2_X4 U2177 ( .A1(n2237), .A2(n2236), .ZN(n2371) );
  INV_X32 U2178 ( .A(x[2]), .ZN(net155744) );
  NAND2_X2 U2179 ( .A1(n2353), .A2(n519), .ZN(net154905) );
  INV_X4 U2180 ( .A(n2718), .ZN(n2650) );
  INV_X4 U2181 ( .A(n1408), .ZN(n1327) );
  NOR2_X4 U2182 ( .A1(net156181), .A2(n729), .ZN(net154290) );
  INV_X4 U2183 ( .A(n1094), .ZN(n2132) );
  NAND2_X4 U2184 ( .A1(net154682), .A2(net154742), .ZN(n2364) );
  NAND2_X4 U2185 ( .A1(n1056), .A2(n1057), .ZN(n1059) );
  XNOR2_X1 U2186 ( .A(n1256), .B(n1255), .ZN(n1309) );
  XNOR2_X2 U2187 ( .A(n2366), .B(n2367), .ZN(net154205) );
  XNOR2_X1 U2188 ( .A(n1311), .B(n1310), .ZN(n1312) );
  NAND2_X4 U2189 ( .A1(n970), .A2(n971), .ZN(n972) );
  INV_X4 U2190 ( .A(n1836), .ZN(n971) );
  NAND2_X4 U2191 ( .A1(n1659), .A2(n1619), .ZN(n1652) );
  NAND3_X1 U2192 ( .A1(n2329), .A2(n2330), .A3(n2549), .ZN(n2313) );
  NAND3_X2 U2193 ( .A1(net154956), .A2(n1947), .A3(n1916), .ZN(n1917) );
  NAND3_X2 U2194 ( .A1(n2588), .A2(net153930), .A3(n861), .ZN(n2590) );
  INV_X2 U2195 ( .A(n2364), .ZN(n973) );
  OAI21_X2 U2196 ( .B1(n1486), .B2(n862), .A(n1485), .ZN(n1699) );
  OAI21_X1 U2197 ( .B1(n1148), .B2(net155827), .A(n1386), .ZN(n1527) );
  NAND2_X4 U2198 ( .A1(net154773), .A2(n1112), .ZN(n2166) );
  NAND2_X2 U2199 ( .A1(n1828), .A2(n825), .ZN(n1873) );
  NAND2_X4 U2200 ( .A1(n2621), .A2(n2622), .ZN(n2623) );
  NOR2_X2 U2201 ( .A1(n2596), .A2(n2600), .ZN(n2229) );
  NAND3_X1 U2202 ( .A1(n2797), .A2(n2786), .A3(n2909), .ZN(n2787) );
  NAND2_X4 U2203 ( .A1(n977), .A2(n976), .ZN(n1880) );
  INV_X1 U2204 ( .A(n1871), .ZN(n978) );
  NAND2_X2 U2205 ( .A1(n1225), .A2(n810), .ZN(n979) );
  NAND2_X4 U2206 ( .A1(n941), .A2(n700), .ZN(n980) );
  NAND2_X4 U2207 ( .A1(n979), .A2(n980), .ZN(n1273) );
  INV_X8 U2208 ( .A(n2629), .ZN(n2548) );
  NAND2_X4 U2209 ( .A1(n1437), .A2(n981), .ZN(n983) );
  INV_X4 U2210 ( .A(n1576), .ZN(n981) );
  NAND2_X2 U2211 ( .A1(n984), .A2(n985), .ZN(n987) );
  NAND2_X4 U2212 ( .A1(n986), .A2(n987), .ZN(n1649) );
  INV_X1 U2213 ( .A(n1611), .ZN(n985) );
  NAND2_X2 U2214 ( .A1(n990), .A2(n991), .ZN(result[33]) );
  INV_X4 U2215 ( .A(n2760), .ZN(n988) );
  INV_X1 U2216 ( .A(n588), .ZN(n989) );
  NOR2_X2 U2217 ( .A1(net153617), .A2(n2814), .ZN(n2823) );
  NAND2_X2 U2218 ( .A1(n2893), .A2(n2793), .ZN(n2796) );
  NAND2_X4 U2219 ( .A1(n1067), .A2(n1068), .ZN(n1070) );
  NAND2_X4 U2220 ( .A1(n1065), .A2(n1066), .ZN(n2582) );
  NAND4_X2 U2221 ( .A1(n1052), .A2(n2851), .A3(n2849), .A4(n2848), .ZN(n2853)
         );
  NAND2_X2 U2222 ( .A1(n1393), .A2(n688), .ZN(n1143) );
  INV_X4 U2223 ( .A(n1393), .ZN(n1142) );
  NAND2_X4 U2224 ( .A1(n1373), .A2(n994), .ZN(n1374) );
  NAND2_X2 U2225 ( .A1(n2152), .A2(n2164), .ZN(n1046) );
  NAND2_X4 U2226 ( .A1(n937), .A2(n2514), .ZN(n2350) );
  INV_X32 U2227 ( .A(n1173), .ZN(n2606) );
  INV_X16 U2228 ( .A(n1172), .ZN(n1173) );
  INV_X2 U2229 ( .A(n1421), .ZN(n992) );
  NAND2_X1 U2230 ( .A1(n576), .A2(n606), .ZN(n2450) );
  OAI21_X2 U2231 ( .B1(n2024), .B2(n2025), .A(n2027), .ZN(n1821) );
  OAI21_X2 U2232 ( .B1(n1165), .B2(n1934), .A(n580), .ZN(n1951) );
  AOI211_X4 U2233 ( .C1(n2657), .C2(n828), .A(n2655), .B(n2654), .ZN(n2671) );
  NAND2_X4 U2234 ( .A1(n2817), .A2(net153611), .ZN(n2818) );
  NAND2_X4 U2235 ( .A1(n1901), .A2(n738), .ZN(n1139) );
  NAND2_X4 U2236 ( .A1(n1896), .A2(n1895), .ZN(n1897) );
  NAND2_X1 U2237 ( .A1(n1304), .A2(net155667), .ZN(n1321) );
  NOR2_X2 U2238 ( .A1(net154031), .A2(n838), .ZN(n2096) );
  INV_X8 U2239 ( .A(n2349), .ZN(n2418) );
  BUF_X4 U2240 ( .A(n2789), .Z(n1060) );
  INV_X8 U2241 ( .A(n1884), .ZN(n2342) );
  NAND2_X4 U2242 ( .A1(n1883), .A2(n1895), .ZN(n1884) );
  NAND2_X2 U2243 ( .A1(n996), .A2(n1230), .ZN(n997) );
  NAND2_X2 U2244 ( .A1(n995), .A2(n1224), .ZN(n998) );
  INV_X4 U2245 ( .A(n1230), .ZN(n995) );
  INV_X1 U2246 ( .A(n995), .ZN(n999) );
  INV_X2 U2247 ( .A(net153562), .ZN(net156776) );
  NAND3_X2 U2248 ( .A1(n2783), .A2(n2798), .A3(n2784), .ZN(n2683) );
  NAND2_X4 U2249 ( .A1(n1081), .A2(n2276), .ZN(n2279) );
  NAND2_X2 U2250 ( .A1(net154038), .A2(n730), .ZN(n2150) );
  NAND2_X2 U2251 ( .A1(net154701), .A2(net154700), .ZN(n2003) );
  NAND2_X4 U2252 ( .A1(n2746), .A2(n2695), .ZN(n2841) );
  NAND2_X4 U2253 ( .A1(n1075), .A2(n1076), .ZN(n1078) );
  AOI211_X4 U2254 ( .C1(n2809), .C2(n2767), .A(n2766), .B(n2765), .ZN(n2774)
         );
  INV_X8 U2255 ( .A(n1453), .ZN(n1553) );
  INV_X8 U2256 ( .A(n1406), .ZN(n1307) );
  NAND2_X4 U2257 ( .A1(n1415), .A2(n1416), .ZN(n1149) );
  INV_X16 U2258 ( .A(n1168), .ZN(n1169) );
  NOR3_X4 U2259 ( .A1(n1868), .A2(n801), .A3(n1866), .ZN(n1869) );
  INV_X8 U2260 ( .A(n1102), .ZN(n1118) );
  NAND2_X4 U2261 ( .A1(n1285), .A2(net155873), .ZN(n1292) );
  NAND2_X4 U2262 ( .A1(n1417), .A2(n1240), .ZN(n1241) );
  NAND2_X2 U2263 ( .A1(n1245), .A2(n1219), .ZN(n1246) );
  NAND3_X4 U2264 ( .A1(net154481), .A2(n2224), .A3(n2223), .ZN(n1002) );
  NAND3_X2 U2265 ( .A1(net154481), .A2(n2224), .A3(n2223), .ZN(n2559) );
  XNOR2_X2 U2266 ( .A(n2564), .B(n2563), .ZN(net154143) );
  NAND2_X4 U2267 ( .A1(n2568), .A2(n509), .ZN(net153701) );
  NAND2_X4 U2268 ( .A1(n2143), .A2(n2142), .ZN(n2144) );
  INV_X8 U2269 ( .A(n1411), .ZN(n1475) );
  NAND2_X4 U2270 ( .A1(n1729), .A2(n1728), .ZN(n2337) );
  NAND2_X4 U2271 ( .A1(n1946), .A2(n1945), .ZN(n1914) );
  OAI21_X4 U2272 ( .B1(n1098), .B2(n2593), .A(net153672), .ZN(n2645) );
  NAND2_X4 U2273 ( .A1(net156482), .A2(net153829), .ZN(net154180) );
  NAND2_X4 U2274 ( .A1(n584), .A2(n2270), .ZN(n2172) );
  NAND2_X2 U2275 ( .A1(n1687), .A2(n1593), .ZN(n1007) );
  NAND2_X4 U2276 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NAND2_X4 U2277 ( .A1(n1007), .A2(n1008), .ZN(n1648) );
  INV_X4 U2278 ( .A(n1593), .ZN(n1006) );
  OAI21_X2 U2279 ( .B1(n2710), .B2(n2800), .A(n2709), .ZN(n2711) );
  OAI21_X2 U2280 ( .B1(n2800), .B2(n2799), .A(n2798), .ZN(n2801) );
  XNOR2_X2 U2281 ( .A(n2647), .B(n2646), .ZN(n2764) );
  NAND3_X4 U2282 ( .A1(n2348), .A2(net156131), .A3(n2524), .ZN(n2349) );
  INV_X8 U2283 ( .A(n1993), .ZN(n1952) );
  NAND2_X4 U2284 ( .A1(n1101), .A2(n1100), .ZN(n1765) );
  INV_X8 U2285 ( .A(n1992), .ZN(n2340) );
  AOI22_X4 U2286 ( .A1(net154155), .A2(n2428), .B1(n622), .B2(n2428), .ZN(
        n2434) );
  NAND2_X4 U2287 ( .A1(n529), .A2(n2386), .ZN(n2661) );
  INV_X2 U2288 ( .A(n1512), .ZN(n1515) );
  INV_X1 U2289 ( .A(n1511), .ZN(n1509) );
  OAI21_X2 U2290 ( .B1(n1751), .B2(n1750), .A(n1749), .ZN(n1887) );
  NAND2_X2 U2291 ( .A1(n2245), .A2(n2244), .ZN(n2246) );
  INV_X8 U2292 ( .A(n2506), .ZN(n1168) );
  INV_X8 U2293 ( .A(n1850), .ZN(n1013) );
  INV_X1 U2294 ( .A(n958), .ZN(n1014) );
  INV_X2 U2295 ( .A(n1014), .ZN(n1015) );
  NAND2_X1 U2296 ( .A1(n2629), .A2(n617), .ZN(n2311) );
  XNOR2_X1 U2297 ( .A(n2579), .B(n2578), .ZN(n2416) );
  INV_X2 U2298 ( .A(n1049), .ZN(n2221) );
  OAI21_X2 U2299 ( .B1(n1871), .B2(n1870), .A(n502), .ZN(n1820) );
  AOI21_X4 U2300 ( .B1(n2089), .B2(n2465), .A(n2376), .ZN(n1016) );
  NAND2_X4 U2301 ( .A1(n2777), .A2(n2776), .ZN(n1017) );
  NAND2_X4 U2302 ( .A1(n1078), .A2(n1077), .ZN(n2777) );
  NAND2_X2 U2303 ( .A1(n2071), .A2(net156803), .ZN(n1019) );
  NAND2_X4 U2304 ( .A1(n1018), .A2(net157076), .ZN(n1020) );
  NAND2_X4 U2305 ( .A1(n1019), .A2(n1020), .ZN(n2569) );
  INV_X4 U2306 ( .A(n2071), .ZN(n1018) );
  INV_X1 U2307 ( .A(net156181), .ZN(net157076) );
  OAI21_X2 U2308 ( .B1(n2070), .B2(n2069), .A(n2068), .ZN(n2071) );
  NAND2_X4 U2309 ( .A1(n509), .A2(n2159), .ZN(n2103) );
  NAND2_X4 U2310 ( .A1(n2568), .A2(n2569), .ZN(n2177) );
  INV_X2 U2311 ( .A(n2569), .ZN(n2309) );
  INV_X4 U2312 ( .A(n2265), .ZN(n2762) );
  XNOR2_X2 U2313 ( .A(n749), .B(n1021), .ZN(n2660) );
  OAI22_X4 U2314 ( .A1(n1174), .A2(n2362), .B1(net155869), .B2(n2472), .ZN(
        n2366) );
  NAND2_X2 U2315 ( .A1(n2475), .A2(n2474), .ZN(n1025) );
  NAND2_X4 U2316 ( .A1(n1023), .A2(n1024), .ZN(n1026) );
  NAND2_X4 U2317 ( .A1(n1025), .A2(n1026), .ZN(n2864) );
  INV_X4 U2318 ( .A(n2475), .ZN(n1023) );
  INV_X4 U2319 ( .A(n2474), .ZN(n1024) );
  NOR2_X2 U2320 ( .A1(n2864), .A2(n2730), .ZN(n2734) );
  INV_X8 U2321 ( .A(n2864), .ZN(n2584) );
  NAND2_X4 U2322 ( .A1(n2330), .A2(n2329), .ZN(net154332) );
  NAND2_X4 U2323 ( .A1(n914), .A2(n592), .ZN(n1561) );
  INV_X2 U2324 ( .A(n2655), .ZN(n2643) );
  NAND2_X4 U2325 ( .A1(n1903), .A2(n1902), .ZN(n1027) );
  NAND2_X2 U2326 ( .A1(n1030), .A2(net157038), .ZN(n1032) );
  NAND2_X4 U2327 ( .A1(n1031), .A2(n1032), .ZN(n2878) );
  XNOR2_X2 U2328 ( .A(n2544), .B(n2878), .ZN(result[30]) );
  NOR2_X4 U2329 ( .A1(n2677), .A2(n2678), .ZN(n2680) );
  NAND2_X4 U2330 ( .A1(n2359), .A2(n2361), .ZN(n2399) );
  NAND2_X2 U2331 ( .A1(n2750), .A2(n2703), .ZN(n1035) );
  NAND2_X2 U2332 ( .A1(n1036), .A2(n1035), .ZN(result[32]) );
  INV_X2 U2333 ( .A(n2750), .ZN(n1033) );
  NAND2_X4 U2334 ( .A1(n1038), .A2(n1039), .ZN(n1041) );
  NAND2_X4 U2335 ( .A1(n1040), .A2(n1041), .ZN(n2387) );
  NAND2_X4 U2336 ( .A1(n2387), .A2(n2386), .ZN(n2511) );
  INV_X2 U2337 ( .A(n2863), .ZN(n2865) );
  NAND2_X4 U2338 ( .A1(n2398), .A2(n2397), .ZN(n2579) );
  NOR2_X2 U2339 ( .A1(n2480), .A2(net154091), .ZN(n2481) );
  NAND2_X4 U2340 ( .A1(net155482), .A2(net155511), .ZN(n1042) );
  XNOR2_X2 U2341 ( .A(n1043), .B(n1914), .ZN(n2336) );
  NAND3_X2 U2342 ( .A1(net154731), .A2(net154728), .A3(net154630), .ZN(
        net154795) );
  NAND2_X4 U2343 ( .A1(net154796), .A2(net154795), .ZN(n2093) );
  XNOR2_X1 U2344 ( .A(n1185), .B(n1189), .ZN(result[1]) );
  NAND2_X4 U2345 ( .A1(n1044), .A2(n1045), .ZN(n1047) );
  NAND2_X4 U2346 ( .A1(n1046), .A2(n1047), .ZN(n2324) );
  INV_X2 U2347 ( .A(n2152), .ZN(n1044) );
  INV_X4 U2348 ( .A(n2164), .ZN(n1045) );
  INV_X4 U2349 ( .A(n2219), .ZN(n1048) );
  INV_X8 U2350 ( .A(n1048), .ZN(n1049) );
  INV_X4 U2351 ( .A(n2549), .ZN(n2550) );
  NAND2_X4 U2352 ( .A1(n1895), .A2(n897), .ZN(n1993) );
  NAND2_X2 U2353 ( .A1(n1807), .A2(n1812), .ZN(n1592) );
  NAND2_X4 U2354 ( .A1(n2513), .A2(n2512), .ZN(n2813) );
  INV_X4 U2355 ( .A(n2114), .ZN(n1154) );
  INV_X8 U2356 ( .A(n2146), .ZN(n2163) );
  INV_X8 U2357 ( .A(n2551), .ZN(n2558) );
  AOI21_X4 U2358 ( .B1(n2434), .B2(n2433), .A(n2432), .ZN(n2435) );
  XNOR2_X1 U2359 ( .A(net154694), .B(net154721), .ZN(n2135) );
  NAND2_X4 U2360 ( .A1(n697), .A2(n1371), .ZN(n1372) );
  NAND2_X4 U2361 ( .A1(x[4]), .A2(n2606), .ZN(n1250) );
  INV_X4 U2362 ( .A(n2128), .ZN(n2129) );
  NAND2_X4 U2363 ( .A1(n1164), .A2(n1163), .ZN(n2555) );
  NOR2_X4 U2364 ( .A1(x[2]), .A2(x[1]), .ZN(n1051) );
  NAND2_X4 U2365 ( .A1(n2408), .A2(n2240), .ZN(n2216) );
  NAND2_X4 U2366 ( .A1(n1233), .A2(n1234), .ZN(n1264) );
  NAND3_X2 U2367 ( .A1(n2894), .A2(n2898), .A3(n2895), .ZN(n1052) );
  INV_X4 U2368 ( .A(n2534), .ZN(n1054) );
  NAND2_X2 U2369 ( .A1(n1058), .A2(n1059), .ZN(n2856) );
  INV_X4 U2370 ( .A(n2855), .ZN(n1057) );
  NAND2_X4 U2371 ( .A1(n2788), .A2(n2787), .ZN(n2898) );
  INV_X2 U2372 ( .A(n2845), .ZN(n2905) );
  NAND2_X4 U2373 ( .A1(n846), .A2(n2535), .ZN(n2614) );
  INV_X1 U2374 ( .A(n1883), .ZN(n1061) );
  NAND2_X1 U2375 ( .A1(n1564), .A2(n1565), .ZN(n1062) );
  NAND2_X2 U2376 ( .A1(n1565), .A2(n1564), .ZN(n1603) );
  NAND2_X4 U2377 ( .A1(n715), .A2(n2115), .ZN(n2202) );
  NOR3_X2 U2378 ( .A1(n1990), .A2(n2342), .A3(n1989), .ZN(n2218) );
  NAND2_X4 U2379 ( .A1(n1063), .A2(n1064), .ZN(n1066) );
  NAND2_X1 U2380 ( .A1(n2443), .A2(n809), .ZN(n1069) );
  INV_X1 U2381 ( .A(n809), .ZN(n1068) );
  INV_X16 U2382 ( .A(n1166), .ZN(n1167) );
  OAI21_X4 U2383 ( .B1(n795), .B2(n2696), .A(n549), .ZN(n2699) );
  OAI21_X2 U2384 ( .B1(n1874), .B2(n1873), .A(n1872), .ZN(n1875) );
  NAND2_X2 U2385 ( .A1(n2879), .A2(n2878), .ZN(n2836) );
  XNOR2_X1 U2386 ( .A(n548), .B(n564), .ZN(n1389) );
  NAND2_X4 U2387 ( .A1(n2592), .A2(net153633), .ZN(net153672) );
  XNOR2_X1 U2388 ( .A(n1958), .B(net157139), .ZN(n1949) );
  NAND2_X4 U2389 ( .A1(n1072), .A2(net156869), .ZN(n1074) );
  NAND2_X4 U2390 ( .A1(n1074), .A2(n1073), .ZN(n1081) );
  INV_X8 U2391 ( .A(n1349), .ZN(n1518) );
  INV_X4 U2392 ( .A(n2483), .ZN(n2487) );
  NAND2_X2 U2393 ( .A1(n2775), .A2(n2900), .ZN(n1077) );
  INV_X4 U2394 ( .A(n2900), .ZN(n1075) );
  NAND2_X4 U2395 ( .A1(n854), .A2(n2876), .ZN(n2778) );
  INV_X2 U2396 ( .A(n1642), .ZN(n1646) );
  XNOR2_X2 U2397 ( .A(n2620), .B(n2652), .ZN(n1080) );
  NAND3_X4 U2398 ( .A1(n1304), .A2(net155667), .A3(net155777), .ZN(n1249) );
  NAND2_X2 U2399 ( .A1(n1092), .A2(n1493), .ZN(n1355) );
  NAND2_X4 U2400 ( .A1(net154334), .A2(n2511), .ZN(net154477) );
  OAI221_X4 U2401 ( .B1(n1169), .B2(n698), .C1(n2225), .C2(net154479), .A(
        net154480), .ZN(n2564) );
  OAI211_X4 U2402 ( .C1(n1412), .C2(n673), .A(n508), .B(n1475), .ZN(n1423) );
  NAND2_X4 U2403 ( .A1(n1287), .A2(n1286), .ZN(n1226) );
  NAND2_X2 U2404 ( .A1(n2508), .A2(net154055), .ZN(n2517) );
  INV_X4 U2405 ( .A(net153875), .ZN(net153876) );
  NAND2_X2 U2406 ( .A1(n2631), .A2(net153875), .ZN(n2385) );
  NAND3_X1 U2407 ( .A1(n1280), .A2(n1335), .A3(n1333), .ZN(n1337) );
  NAND3_X2 U2408 ( .A1(net158266), .A2(n2808), .A3(n2807), .ZN(n2810) );
  NAND3_X2 U2409 ( .A1(net153633), .A2(n2806), .A3(n2805), .ZN(net153630) );
  NAND2_X2 U2410 ( .A1(n2805), .A2(n2806), .ZN(n2543) );
  NAND2_X4 U2411 ( .A1(n1170), .A2(net156089), .ZN(n2667) );
  NAND2_X4 U2412 ( .A1(n2791), .A2(n2792), .ZN(n2793) );
  NAND3_X2 U2413 ( .A1(n2665), .A2(n833), .A3(n2658), .ZN(net156810) );
  INV_X4 U2414 ( .A(net156810), .ZN(net156811) );
  XNOR2_X1 U2415 ( .A(n848), .B(n1269), .ZN(result[4]) );
  XNOR2_X1 U2416 ( .A(n1984), .B(n596), .ZN(result[20]) );
  AOI21_X1 U2417 ( .B1(n596), .B2(n1988), .A(n1987), .ZN(n2015) );
  NAND2_X1 U2418 ( .A1(n596), .A2(n2166), .ZN(n2173) );
  AOI22_X2 U2419 ( .A1(net154423), .A2(n596), .B1(n2567), .B2(n2565), .ZN(
        n2300) );
  XNOR2_X2 U2420 ( .A(n1933), .B(n520), .ZN(n1083) );
  NAND2_X1 U2421 ( .A1(n1079), .A2(n1652), .ZN(n1629) );
  NAND2_X4 U2422 ( .A1(n2163), .A2(n2162), .ZN(n2151) );
  AOI21_X2 U2423 ( .B1(n2182), .B2(net153533), .A(n2181), .ZN(n2183) );
  NAND2_X1 U2424 ( .A1(n2288), .A2(net153533), .ZN(n2180) );
  NAND2_X4 U2425 ( .A1(n2118), .A2(n2119), .ZN(n2390) );
  NAND2_X4 U2426 ( .A1(n1787), .A2(n1297), .ZN(n1598) );
  NOR2_X4 U2427 ( .A1(n1085), .A2(net155985), .ZN(n1084) );
  XNOR2_X2 U2428 ( .A(net154606), .B(net156664), .ZN(n1095) );
  NAND2_X4 U2429 ( .A1(n2253), .A2(n2252), .ZN(n2268) );
  INV_X1 U2430 ( .A(n1650), .ZN(n1086) );
  INV_X32 U2431 ( .A(x[0]), .ZN(net156745) );
  INV_X2 U2432 ( .A(n2099), .ZN(n1087) );
  NAND2_X4 U2433 ( .A1(n1344), .A2(n1345), .ZN(n1315) );
  NAND3_X2 U2434 ( .A1(n1197), .A2(n956), .A3(n1196), .ZN(n1216) );
  NAND2_X4 U2435 ( .A1(n1465), .A2(n1464), .ZN(n1736) );
  OAI21_X1 U2436 ( .B1(n900), .B2(net155835), .A(n2111), .ZN(n2276) );
  OAI21_X1 U2437 ( .B1(n2112), .B2(net155869), .A(n2049), .ZN(n2050) );
  NOR2_X4 U2438 ( .A1(x[13]), .A2(x[14]), .ZN(n1088) );
  NAND2_X4 U2439 ( .A1(n2690), .A2(n2689), .ZN(net153796) );
  INV_X1 U2440 ( .A(n2356), .ZN(n1089) );
  INV_X8 U2441 ( .A(n2646), .ZN(n2653) );
  XNOR2_X2 U2442 ( .A(n2411), .B(n2412), .ZN(n1090) );
  NOR2_X2 U2443 ( .A1(n1910), .A2(n518), .ZN(n1913) );
  INV_X8 U2444 ( .A(n1714), .ZN(n1715) );
  INV_X1 U2445 ( .A(n2431), .ZN(n2398) );
  OAI21_X1 U2446 ( .B1(n821), .B2(net155827), .A(n1982), .ZN(n2270) );
  INV_X4 U2447 ( .A(n2048), .ZN(n2112) );
  NAND2_X1 U2448 ( .A1(n549), .A2(net153532), .ZN(n2421) );
  NAND2_X4 U2449 ( .A1(net158117), .A2(net153621), .ZN(n2516) );
  NOR2_X4 U2450 ( .A1(x[13]), .A2(x[14]), .ZN(n1091) );
  OAI21_X4 U2451 ( .B1(n2617), .B2(n2676), .A(n860), .ZN(n2619) );
  INV_X1 U2452 ( .A(n1783), .ZN(n1711) );
  OAI22_X4 U2453 ( .A1(net155885), .A2(n2461), .B1(n2594), .B2(net155857), 
        .ZN(n2535) );
  OAI21_X4 U2454 ( .B1(n1346), .B2(n1347), .A(n1363), .ZN(n1092) );
  OAI221_X4 U2455 ( .B1(n1838), .B2(n1912), .C1(n513), .C2(n600), .A(n607), 
        .ZN(n1901) );
  NAND2_X4 U2456 ( .A1(n1600), .A2(n1599), .ZN(n1714) );
  NOR2_X4 U2457 ( .A1(n1598), .A2(n956), .ZN(n1599) );
  NAND3_X2 U2458 ( .A1(net154629), .A2(net154630), .A3(n2055), .ZN(n1093) );
  NAND3_X2 U2459 ( .A1(net154630), .A2(net154629), .A3(n2055), .ZN(n2596) );
  INV_X2 U2460 ( .A(n1519), .ZN(n1358) );
  NAND2_X4 U2461 ( .A1(net154742), .A2(n2046), .ZN(n1094) );
  NAND2_X4 U2462 ( .A1(n1718), .A2(net156073), .ZN(n1745) );
  NAND2_X4 U2463 ( .A1(net154616), .A2(n2129), .ZN(n2131) );
  NAND2_X4 U2464 ( .A1(n2141), .A2(n2140), .ZN(net153613) );
  NAND2_X4 U2465 ( .A1(n2458), .A2(n2611), .ZN(n2539) );
  NAND2_X4 U2466 ( .A1(n1096), .A2(n1097), .ZN(net154578) );
  NAND2_X4 U2467 ( .A1(n2279), .A2(n2278), .ZN(n2280) );
  NOR3_X4 U2468 ( .A1(n2699), .A2(n2697), .A3(n2698), .ZN(net153674) );
  INV_X4 U2469 ( .A(net154291), .ZN(net154602) );
  NAND4_X4 U2470 ( .A1(n1810), .A2(n1809), .A3(n1808), .A4(n1807), .ZN(n1811)
         );
  NAND3_X2 U2471 ( .A1(n1539), .A2(n1540), .A3(n1541), .ZN(n1636) );
  INV_X4 U2472 ( .A(n1540), .ZN(n1619) );
  NAND2_X4 U2473 ( .A1(n2755), .A2(n2756), .ZN(n2757) );
  NAND2_X4 U2474 ( .A1(n2754), .A2(n2753), .ZN(n2755) );
  NOR2_X2 U2475 ( .A1(n2339), .A2(n2340), .ZN(n2344) );
  NOR3_X2 U2476 ( .A1(n2243), .A2(n2242), .A3(n2241), .ZN(n2245) );
  NAND2_X4 U2477 ( .A1(n1790), .A2(n1789), .ZN(n1102) );
  INV_X8 U2478 ( .A(n1135), .ZN(n1789) );
  INV_X8 U2479 ( .A(n2274), .ZN(n2306) );
  INV_X4 U2480 ( .A(n1324), .ZN(n1298) );
  INV_X8 U2481 ( .A(n1662), .ZN(n1741) );
  NAND2_X1 U2482 ( .A1(n1409), .A2(n1327), .ZN(n1106) );
  NAND2_X2 U2483 ( .A1(n1104), .A2(n1105), .ZN(n1107) );
  NAND2_X4 U2484 ( .A1(n1106), .A2(n1107), .ZN(n1380) );
  INV_X1 U2485 ( .A(n1409), .ZN(n1104) );
  INV_X4 U2486 ( .A(n1327), .ZN(n1105) );
  NAND2_X2 U2487 ( .A1(n1325), .A2(n516), .ZN(n1109) );
  NAND2_X4 U2488 ( .A1(n1108), .A2(net155482), .ZN(n1110) );
  NAND2_X4 U2489 ( .A1(n1109), .A2(n1110), .ZN(n1381) );
  INV_X4 U2490 ( .A(n1325), .ZN(n1108) );
  NAND2_X2 U2491 ( .A1(n1380), .A2(n1407), .ZN(n1383) );
  XNOR2_X1 U2492 ( .A(n1274), .B(n1273), .ZN(n1276) );
  XNOR2_X1 U2493 ( .A(n2492), .B(n1167), .ZN(n1111) );
  INV_X2 U2494 ( .A(n1963), .ZN(n1112) );
  NAND2_X2 U2495 ( .A1(net155496), .A2(n1418), .ZN(n1114) );
  NAND2_X4 U2496 ( .A1(n1113), .A2(x[9]), .ZN(n1115) );
  NAND2_X4 U2497 ( .A1(n1114), .A2(n1115), .ZN(n1575) );
  NOR2_X2 U2498 ( .A1(n1152), .A2(n1039), .ZN(n2233) );
  INV_X4 U2499 ( .A(n1017), .ZN(n2857) );
  NAND3_X4 U2500 ( .A1(n1211), .A2(n1210), .A3(n1212), .ZN(net155697) );
  NAND2_X4 U2501 ( .A1(n1209), .A2(n1051), .ZN(n1212) );
  AOI22_X4 U2502 ( .A1(x[2]), .A2(x[3]), .B1(x[1]), .B2(x[3]), .ZN(n1211) );
  OAI21_X4 U2503 ( .B1(n642), .B2(n2128), .A(n2130), .ZN(n2086) );
  NAND3_X4 U2504 ( .A1(net155775), .A2(net155744), .A3(net155508), .ZN(n1116)
         );
  NAND3_X4 U2505 ( .A1(net155775), .A2(net155744), .A3(net155508), .ZN(n1117)
         );
  OAI21_X2 U2506 ( .B1(n2338), .B2(n822), .A(n2337), .ZN(n2339) );
  NAND2_X2 U2507 ( .A1(n593), .A2(n577), .ZN(n1482) );
  NAND2_X4 U2508 ( .A1(n2790), .A2(n2851), .ZN(n2792) );
  OAI22_X4 U2509 ( .A1(n1175), .A2(n2461), .B1(net155869), .B2(n2594), .ZN(
        n2459) );
  OAI21_X1 U2510 ( .B1(net155827), .B2(n2472), .A(n2471), .ZN(n2581) );
  NAND2_X4 U2511 ( .A1(n2809), .A2(n2651), .ZN(n2848) );
  OAI22_X4 U2512 ( .A1(n1174), .A2(n2361), .B1(net155869), .B2(n2542), .ZN(
        n2405) );
  NAND2_X4 U2513 ( .A1(n2360), .A2(n2399), .ZN(n2542) );
  NAND4_X2 U2514 ( .A1(n2344), .A2(net153613), .A3(n2343), .A4(net154293), 
        .ZN(n2419) );
  OAI21_X4 U2515 ( .B1(n2859), .B2(n2882), .A(n2858), .ZN(n2861) );
  NOR2_X4 U2516 ( .A1(n2844), .A2(n2843), .ZN(n2859) );
  NAND2_X4 U2517 ( .A1(net153700), .A2(n553), .ZN(n2298) );
  NAND3_X2 U2518 ( .A1(n695), .A2(n2284), .A3(n2285), .ZN(n2294) );
  OAI21_X2 U2519 ( .B1(n1148), .B2(net155869), .A(n1285), .ZN(n1284) );
  NAND2_X4 U2520 ( .A1(n1270), .A2(n1271), .ZN(n1272) );
  AOI21_X4 U2521 ( .B1(n1524), .B2(n1523), .A(n1522), .ZN(n1532) );
  NOR2_X4 U2522 ( .A1(n1138), .A2(n2267), .ZN(n2299) );
  INV_X4 U2523 ( .A(n2216), .ZN(n2209) );
  NOR2_X2 U2524 ( .A1(n1677), .A2(n1171), .ZN(n1679) );
  NAND2_X4 U2525 ( .A1(n1139), .A2(n1140), .ZN(n1903) );
  NAND2_X2 U2526 ( .A1(n2680), .A2(n2609), .ZN(n2785) );
  NAND2_X4 U2527 ( .A1(n1880), .A2(n1879), .ZN(n1992) );
  NOR2_X4 U2528 ( .A1(n2347), .A2(n2346), .ZN(n2348) );
  NAND2_X4 U2529 ( .A1(n1119), .A2(n1120), .ZN(n1122) );
  NAND2_X2 U2530 ( .A1(n1122), .A2(n1121), .ZN(result[35]) );
  INV_X4 U2531 ( .A(n2918), .ZN(n1119) );
  INV_X4 U2532 ( .A(n2917), .ZN(n1120) );
  INV_X8 U2533 ( .A(n1725), .ZN(n1871) );
  OAI21_X2 U2534 ( .B1(n1956), .B2(n1774), .A(n1773), .ZN(n1826) );
  NAND2_X4 U2535 ( .A1(n1895), .A2(n1883), .ZN(n1125) );
  NAND2_X4 U2536 ( .A1(n1128), .A2(n1129), .ZN(n1829) );
  OAI21_X1 U2537 ( .B1(net155827), .B2(n2686), .A(n2685), .ZN(n2830) );
  OAI21_X1 U2538 ( .B1(net155839), .B2(n545), .A(n2595), .ZN(n2657) );
  NAND2_X2 U2539 ( .A1(net155884), .A2(x[9]), .ZN(n1130) );
  NAND2_X4 U2540 ( .A1(n1456), .A2(n1130), .ZN(n1657) );
  NAND2_X2 U2541 ( .A1(n1569), .A2(n1580), .ZN(n1132) );
  NAND2_X4 U2542 ( .A1(n1131), .A2(n839), .ZN(n1133) );
  NAND2_X4 U2543 ( .A1(n1133), .A2(n1132), .ZN(n1462) );
  XNOR2_X2 U2544 ( .A(n1658), .B(n839), .ZN(n1661) );
  INV_X8 U2545 ( .A(n1581), .ZN(n1569) );
  XNOR2_X2 U2546 ( .A(n1463), .B(n814), .ZN(n1465) );
  NAND2_X4 U2547 ( .A1(n2491), .A2(n2490), .ZN(n2492) );
  OAI22_X1 U2548 ( .A1(n2705), .A2(n1848), .B1(net155827), .B2(n1847), .ZN(
        n1876) );
  OAI21_X2 U2549 ( .B1(net155839), .B2(n1847), .A(n1775), .ZN(n1879) );
  INV_X4 U2550 ( .A(n2363), .ZN(n2208) );
  AOI21_X2 U2551 ( .B1(n1973), .B2(n824), .A(n1971), .ZN(n1974) );
  NAND2_X4 U2552 ( .A1(n1922), .A2(n1921), .ZN(net154858) );
  OAI21_X4 U2553 ( .B1(net156405), .B2(net154856), .A(x[20]), .ZN(net154796)
         );
  INV_X4 U2554 ( .A(n2320), .ZN(n2267) );
  INV_X4 U2555 ( .A(n1779), .ZN(n1780) );
  NAND2_X4 U2556 ( .A1(n2384), .A2(net154234), .ZN(n2499) );
  XNOR2_X1 U2557 ( .A(n2372), .B(n708), .ZN(n2196) );
  NAND2_X1 U2558 ( .A1(n2372), .A2(n2371), .ZN(n2247) );
  NAND2_X1 U2559 ( .A1(n2226), .A2(n2228), .ZN(n2375) );
  NAND2_X1 U2560 ( .A1(n692), .A2(n2228), .ZN(n2125) );
  NAND2_X1 U2561 ( .A1(net156073), .A2(n2228), .ZN(n2193) );
  OAI21_X2 U2562 ( .B1(x[25]), .B2(n2228), .A(x[26]), .ZN(n2230) );
  INV_X8 U2563 ( .A(n1381), .ZN(n1326) );
  NOR2_X4 U2564 ( .A1(n1747), .A2(n530), .ZN(n1134) );
  NAND2_X4 U2565 ( .A1(n1788), .A2(n1088), .ZN(n1135) );
  INV_X1 U2566 ( .A(n2567), .ZN(n1136) );
  INV_X8 U2567 ( .A(n2177), .ZN(n2567) );
  NAND2_X4 U2568 ( .A1(n2500), .A2(n583), .ZN(n2808) );
  NAND2_X4 U2569 ( .A1(n1654), .A2(n1653), .ZN(n1730) );
  NAND2_X4 U2570 ( .A1(n2327), .A2(n2326), .ZN(net153532) );
  OAI211_X4 U2571 ( .C1(n1645), .C2(n1646), .A(n1643), .B(n1644), .ZN(n1725)
         );
  NAND2_X4 U2572 ( .A1(n1142), .A2(n1475), .ZN(n1144) );
  NAND2_X4 U2573 ( .A1(n1143), .A2(n1144), .ZN(n1395) );
  NAND2_X4 U2574 ( .A1(n1525), .A2(n1678), .ZN(n1670) );
  NAND2_X4 U2575 ( .A1(x[4]), .A2(n1212), .ZN(n1304) );
  NAND2_X4 U2576 ( .A1(n2283), .A2(n2282), .ZN(n1985) );
  INV_X2 U2577 ( .A(n1145), .ZN(n1146) );
  NAND2_X2 U2578 ( .A1(n2085), .A2(net154682), .ZN(n2118) );
  INV_X1 U2579 ( .A(n1759), .ZN(n1817) );
  INV_X4 U2580 ( .A(n1603), .ZN(n1566) );
  OAI21_X2 U2581 ( .B1(n2829), .B2(n2828), .A(n2830), .ZN(n2832) );
  NAND2_X4 U2582 ( .A1(n1375), .A2(n1374), .ZN(n1399) );
  NAND2_X4 U2583 ( .A1(n1666), .A2(n1424), .ZN(n1434) );
  NAND2_X4 U2584 ( .A1(n2258), .A2(n1165), .ZN(n2259) );
  NAND2_X4 U2585 ( .A1(n1154), .A2(n1153), .ZN(n1156) );
  NAND2_X4 U2586 ( .A1(n1759), .A2(n771), .ZN(n1704) );
  NAND2_X2 U2587 ( .A1(n2821), .A2(n2811), .ZN(n2846) );
  OAI21_X2 U2588 ( .B1(n1626), .B2(n1625), .A(n1642), .ZN(n1627) );
  INV_X4 U2589 ( .A(n1092), .ZN(n1676) );
  INV_X8 U2590 ( .A(n2529), .ZN(n2530) );
  NAND2_X4 U2591 ( .A1(n860), .A2(n2676), .ZN(n2784) );
  NAND2_X4 U2592 ( .A1(n1414), .A2(n994), .ZN(n1415) );
  NAND2_X4 U2593 ( .A1(n1636), .A2(n1071), .ZN(n1594) );
  NAND2_X1 U2594 ( .A1(n1472), .A2(n932), .ZN(n1439) );
  NAND2_X1 U2595 ( .A1(n1571), .A2(n932), .ZN(n1440) );
  NOR2_X4 U2596 ( .A1(net153562), .A2(n2857), .ZN(n2858) );
  NAND2_X4 U2597 ( .A1(n2612), .A2(n2611), .ZN(n2677) );
  NAND2_X4 U2598 ( .A1(n2229), .A2(n2598), .ZN(n2358) );
  OAI21_X2 U2599 ( .B1(net155837), .B2(n1183), .A(net157416), .ZN(n1207) );
  NAND2_X1 U2600 ( .A1(n1215), .A2(n1214), .ZN(n1219) );
  NAND2_X4 U2601 ( .A1(n1315), .A2(n1306), .ZN(n1361) );
  NAND2_X1 U2602 ( .A1(n1807), .A2(n1809), .ZN(n1697) );
  XNOR2_X1 U2603 ( .A(n1623), .B(n1637), .ZN(n1622) );
  NAND2_X4 U2604 ( .A1(n1322), .A2(n1323), .ZN(n1408) );
  NAND2_X4 U2605 ( .A1(n2548), .A2(n1169), .ZN(net154334) );
  INV_X8 U2606 ( .A(net154332), .ZN(net154481) );
  NAND2_X4 U2607 ( .A1(n2374), .A2(n2373), .ZN(net154247) );
  NAND2_X4 U2608 ( .A1(n1800), .A2(n1799), .ZN(n1803) );
  OAI21_X1 U2609 ( .B1(net155827), .B2(n2212), .A(n2211), .ZN(n2552) );
  INV_X4 U2610 ( .A(n2115), .ZN(n1153) );
  NAND3_X2 U2611 ( .A1(n2892), .A2(n2893), .A3(n2772), .ZN(n2724) );
  INV_X8 U2612 ( .A(n2679), .ZN(n2540) );
  NAND2_X4 U2613 ( .A1(n1281), .A2(n943), .ZN(n1282) );
  XNOR2_X1 U2614 ( .A(net156989), .B(net154905), .ZN(n2354) );
  NAND2_X4 U2615 ( .A1(n2717), .A2(n2479), .ZN(n2484) );
  NAND2_X1 U2616 ( .A1(n2841), .A2(net153674), .ZN(n2701) );
  NAND3_X2 U2617 ( .A1(n2248), .A2(n2247), .A3(n2246), .ZN(net154322) );
  NAND2_X4 U2618 ( .A1(n2400), .A2(n2461), .ZN(n2462) );
  NAND2_X4 U2619 ( .A1(n2401), .A2(n2462), .ZN(n2594) );
  INV_X8 U2620 ( .A(n2462), .ZN(n2468) );
  NAND2_X4 U2621 ( .A1(n2619), .A2(n2783), .ZN(n2646) );
  OAI21_X2 U2622 ( .B1(net155839), .B2(n2212), .A(n2126), .ZN(n2658) );
  INV_X8 U2623 ( .A(n1180), .ZN(n1181) );
  OAI21_X1 U2624 ( .B1(net155827), .B2(n2093), .A(n2092), .ZN(n2273) );
  NAND2_X4 U2625 ( .A1(n1795), .A2(n1801), .ZN(n1796) );
  INV_X8 U2626 ( .A(n2835), .ZN(n2882) );
  NAND3_X2 U2627 ( .A1(n2671), .A2(n2769), .A3(n576), .ZN(n2743) );
  INV_X4 U2628 ( .A(n2556), .ZN(n1158) );
  NAND2_X4 U2629 ( .A1(n2762), .A2(n2761), .ZN(n2566) );
  NAND2_X4 U2630 ( .A1(n1284), .A2(n1283), .ZN(n1405) );
  INV_X8 U2631 ( .A(n1575), .ZN(n1596) );
  NAND2_X4 U2632 ( .A1(n1948), .A2(n1969), .ZN(net154285) );
  NAND2_X4 U2633 ( .A1(n1805), .A2(n1806), .ZN(n1968) );
  NAND2_X4 U2634 ( .A1(n1481), .A2(n1480), .ZN(n1695) );
  NOR3_X4 U2635 ( .A1(n1990), .A2(n2342), .A3(n1989), .ZN(n1954) );
  NAND2_X4 U2636 ( .A1(n2833), .A2(n2834), .ZN(n2835) );
  NAND2_X4 U2637 ( .A1(n2806), .A2(n2805), .ZN(net153784) );
  NAND4_X4 U2638 ( .A1(n2670), .A2(n2723), .A3(n2526), .A4(n2527), .ZN(n2806)
         );
  INV_X8 U2639 ( .A(n2113), .ZN(n2130) );
  INV_X32 U2640 ( .A(x[18]), .ZN(net154940) );
  INV_X32 U2641 ( .A(x[17]), .ZN(net154947) );
  NAND2_X1 U2642 ( .A1(n2477), .A2(n549), .ZN(n2317) );
  OAI211_X1 U2643 ( .C1(n1986), .C2(net154760), .A(n587), .B(n1112), .ZN(n1988) );
  NAND2_X4 U2644 ( .A1(net157139), .A2(n2522), .ZN(n2043) );
  NAND2_X4 U2645 ( .A1(n1548), .A2(n1296), .ZN(n1324) );
  NOR2_X2 U2646 ( .A1(n2587), .A2(n2586), .ZN(n2588) );
  INV_X2 U2647 ( .A(n2234), .ZN(n2238) );
  INV_X4 U2648 ( .A(net154700), .ZN(net154744) );
  NAND2_X4 U2649 ( .A1(n1290), .A2(n1218), .ZN(n1288) );
  AOI21_X4 U2650 ( .B1(n2011), .B2(n2049), .A(n2010), .ZN(net154791) );
  NAND3_X2 U2651 ( .A1(n2770), .A2(n852), .A3(n2739), .ZN(n2740) );
  INV_X8 U2652 ( .A(n1170), .ZN(n2479) );
  NOR3_X2 U2653 ( .A1(n2732), .A2(n571), .A3(n2731), .ZN(n2733) );
  NAND2_X4 U2654 ( .A1(n1545), .A2(n1614), .ZN(n1467) );
  NAND2_X4 U2655 ( .A1(n1452), .A2(n1451), .ZN(n1581) );
  NAND2_X2 U2656 ( .A1(n715), .A2(n2115), .ZN(n1155) );
  NAND2_X4 U2657 ( .A1(n1155), .A2(n1156), .ZN(n2199) );
  OAI21_X4 U2658 ( .B1(n2132), .B2(n2131), .A(n2130), .ZN(n2133) );
  NAND2_X4 U2659 ( .A1(n2144), .A2(n2145), .ZN(n2146) );
  OAI21_X2 U2660 ( .B1(net153700), .B2(n2567), .A(n553), .ZN(n2318) );
  OAI21_X2 U2661 ( .B1(n2321), .B2(n2320), .A(n549), .ZN(n2425) );
  NAND2_X4 U2662 ( .A1(n1220), .A2(n1226), .ZN(n1245) );
  OAI21_X4 U2663 ( .B1(n816), .B2(n530), .A(n1746), .ZN(n1810) );
  NAND3_X1 U2664 ( .A1(n2269), .A2(n2270), .A3(n2268), .ZN(n2272) );
  XNOR2_X2 U2665 ( .A(net154642), .B(net154848), .ZN(n1998) );
  NAND2_X4 U2666 ( .A1(n2691), .A2(n2692), .ZN(n2694) );
  XNOR2_X1 U2667 ( .A(n1951), .B(n2290), .ZN(result[19]) );
  NOR2_X1 U2668 ( .A1(n2290), .A2(n2167), .ZN(n2168) );
  NOR3_X2 U2669 ( .A1(n1472), .A2(n1473), .A3(n1571), .ZN(n1469) );
  NAND2_X4 U2670 ( .A1(n1648), .A2(n1647), .ZN(n1663) );
  NAND2_X4 U2671 ( .A1(n1913), .A2(n1912), .ZN(n1945) );
  NAND2_X2 U2672 ( .A1(n2556), .A2(n2557), .ZN(n1159) );
  NAND2_X4 U2673 ( .A1(n1157), .A2(n1158), .ZN(n1160) );
  INV_X4 U2674 ( .A(n2557), .ZN(n1157) );
  NAND2_X4 U2675 ( .A1(n1161), .A2(n1162), .ZN(n1164) );
  INV_X4 U2676 ( .A(n2561), .ZN(n1161) );
  INV_X4 U2677 ( .A(n2553), .ZN(n1162) );
  INV_X2 U2678 ( .A(n2560), .ZN(n2553) );
  OAI22_X4 U2679 ( .A1(n1174), .A2(n2057), .B1(net155869), .B2(n2212), .ZN(
        n2083) );
  NAND2_X2 U2680 ( .A1(x[18]), .A2(n1001), .ZN(n1979) );
  INV_X8 U2681 ( .A(n1083), .ZN(n1165) );
  OAI21_X4 U2682 ( .B1(n1751), .B2(n1911), .A(n1099), .ZN(n1912) );
  NAND2_X1 U2683 ( .A1(net158242), .A2(n2105), .ZN(n2107) );
  NAND2_X4 U2684 ( .A1(n1402), .A2(n1408), .ZN(n1404) );
  NAND2_X2 U2685 ( .A1(net153623), .A2(net157773), .ZN(n2449) );
  AOI22_X4 U2686 ( .A1(n2235), .A2(n2414), .B1(n2235), .B2(net155869), .ZN(
        n2195) );
  NAND2_X1 U2687 ( .A1(net158219), .A2(net157527), .ZN(n2819) );
  NAND2_X4 U2688 ( .A1(n2077), .A2(n560), .ZN(n2329) );
  OAI211_X4 U2689 ( .C1(net155379), .C2(net155696), .A(net155777), .B(n1198), 
        .ZN(n1215) );
  OAI22_X4 U2690 ( .A1(n1175), .A2(n2469), .B1(net155869), .B2(n2686), .ZN(
        n2534) );
  OAI22_X1 U2691 ( .A1(n2705), .A2(n1793), .B1(net155827), .B2(n559), .ZN(
        n1958) );
  NAND2_X4 U2692 ( .A1(n1551), .A2(n1550), .ZN(n1609) );
  INV_X8 U2693 ( .A(n1470), .ZN(n1588) );
  NAND4_X4 U2694 ( .A1(n1405), .A2(n1403), .A3(n1404), .A4(n1406), .ZN(n1470)
         );
  NAND2_X4 U2695 ( .A1(n566), .A2(net156614), .ZN(n1838) );
  NOR2_X4 U2696 ( .A1(net158297), .A2(n2363), .ZN(n2365) );
  NAND3_X2 U2697 ( .A1(n2847), .A2(n2824), .A3(n2846), .ZN(n2825) );
  INV_X1 U2698 ( .A(n2897), .ZN(n2900) );
  XNOR2_X1 U2699 ( .A(n2776), .B(n2897), .ZN(n2727) );
  INV_X16 U2700 ( .A(net155855), .ZN(net156073) );
  NOR2_X4 U2701 ( .A1(n1954), .A2(n1953), .ZN(n1955) );
  XNOR2_X1 U2702 ( .A(n2015), .B(n2032), .ZN(result[21]) );
  NAND2_X4 U2703 ( .A1(net154341), .A2(n2220), .ZN(n2187) );
  INV_X1 U2704 ( .A(n833), .ZN(n2662) );
  OAI21_X2 U2705 ( .B1(n2568), .B2(n2306), .A(n2324), .ZN(n2307) );
  NAND3_X2 U2706 ( .A1(n2289), .A2(n1165), .A3(n1985), .ZN(n2293) );
  INV_X8 U2707 ( .A(n1090), .ZN(n1170) );
  INV_X8 U2708 ( .A(n945), .ZN(n1171) );
  INV_X2 U2709 ( .A(n2879), .ZN(n2880) );
  OAI211_X4 U2710 ( .C1(n2774), .C2(n2773), .A(n2772), .B(n2771), .ZN(n2775)
         );
  NAND4_X4 U2711 ( .A1(n2769), .A2(n852), .A3(n2770), .A4(n2894), .ZN(n2771)
         );
  NAND2_X4 U2712 ( .A1(n1436), .A2(n1435), .ZN(n1660) );
  XNOR2_X1 U2713 ( .A(n1512), .B(n1540), .ZN(n1511) );
  NAND2_X4 U2714 ( .A1(net154699), .A2(n2201), .ZN(n2204) );
  INV_X4 U2715 ( .A(n2841), .ZN(n2844) );
  NAND2_X4 U2716 ( .A1(n2455), .A2(n2454), .ZN(n2679) );
  NAND2_X4 U2717 ( .A1(n2244), .A2(n2239), .ZN(n2113) );
  NAND2_X4 U2718 ( .A1(n1298), .A2(net154943), .ZN(n1370) );
  NAND2_X4 U2719 ( .A1(n1370), .A2(x[8]), .ZN(n1457) );
  XNOR2_X1 U2720 ( .A(n1517), .B(n544), .ZN(result[6]) );
  OAI21_X1 U2721 ( .B1(n1518), .B2(n1517), .A(n1516), .ZN(n1354) );
  INV_X4 U2722 ( .A(n2810), .ZN(n2821) );
  XNOR2_X2 U2723 ( .A(n2476), .B(n2864), .ZN(result[29]) );
  NAND2_X4 U2724 ( .A1(n1342), .A2(n1341), .ZN(n1493) );
  NAND2_X4 U2725 ( .A1(n1367), .A2(n1366), .ZN(n1494) );
  NAND2_X1 U2726 ( .A1(net154629), .A2(n1181), .ZN(net156057) );
  OAI21_X4 U2727 ( .B1(n2862), .B2(n2861), .A(n2860), .ZN(n2889) );
  NAND2_X4 U2728 ( .A1(n1908), .A2(n1909), .ZN(n1946) );
  NAND2_X4 U2729 ( .A1(net157139), .A2(n2352), .ZN(n2077) );
  NAND2_X4 U2730 ( .A1(net155315), .A2(n1608), .ZN(n1179) );
  INV_X8 U2731 ( .A(net157615), .ZN(net155315) );
  NAND2_X4 U2732 ( .A1(n1790), .A2(n1789), .ZN(n1791) );
  NAND2_X4 U2733 ( .A1(n2897), .A2(n2898), .ZN(n2851) );
  NAND2_X4 U2734 ( .A1(net153543), .A2(net153540), .ZN(n2697) );
  NAND2_X4 U2735 ( .A1(n2572), .A2(n2571), .ZN(net153541) );
  NAND2_X4 U2736 ( .A1(n1802), .A2(n857), .ZN(n1830) );
  NAND2_X4 U2737 ( .A1(n1798), .A2(n1797), .ZN(net154810) );
  NAND2_X4 U2738 ( .A1(n944), .A2(n2273), .ZN(n2274) );
  NAND2_X4 U2739 ( .A1(n1731), .A2(n1730), .ZN(n1770) );
  AOI21_X4 U2740 ( .B1(n909), .B2(n1768), .A(n1767), .ZN(n1771) );
  NAND2_X4 U2741 ( .A1(n1478), .A2(n1477), .ZN(n1542) );
  NAND2_X4 U2742 ( .A1(n2641), .A2(n2640), .ZN(n2691) );
  NAND2_X4 U2743 ( .A1(n2626), .A2(n2625), .ZN(net153856) );
  AOI21_X4 U2744 ( .B1(net157295), .B2(net158219), .A(n826), .ZN(n2525) );
  NAND2_X4 U2745 ( .A1(n2503), .A2(n2502), .ZN(n2718) );
  NAND2_X4 U2746 ( .A1(n2856), .A2(n2907), .ZN(net153560) );
  XNOR2_X1 U2747 ( .A(n1460), .B(n834), .ZN(result[10]) );
  NAND2_X4 U2748 ( .A1(n1215), .A2(n1214), .ZN(n1290) );
  INV_X8 U2749 ( .A(n2199), .ZN(n2205) );
  NAND2_X4 U2750 ( .A1(n2365), .A2(n1094), .ZN(n2454) );
  OAI22_X2 U2751 ( .A1(n1676), .A2(n1675), .B1(n1677), .B2(n1171), .ZN(n1495)
         );
  NOR3_X4 U2752 ( .A1(n1786), .A2(n537), .A3(n1785), .ZN(n1792) );
  NAND2_X4 U2753 ( .A1(n2455), .A2(n2454), .ZN(n2609) );
  NOR2_X4 U2754 ( .A1(n2215), .A2(n2216), .ZN(n2217) );
  NAND2_X4 U2755 ( .A1(n1942), .A2(n1943), .ZN(net154879) );
  NAND2_X2 U2756 ( .A1(n2209), .A2(n2214), .ZN(n2210) );
  NAND2_X4 U2757 ( .A1(n1250), .A2(n1249), .ZN(n1256) );
  NAND2_X4 U2758 ( .A1(n1307), .A2(n1280), .ZN(n1377) );
  INV_X8 U2759 ( .A(n863), .ZN(n2074) );
  NAND2_X4 U2760 ( .A1(n1765), .A2(n1891), .ZN(n1878) );
  OAI211_X4 U2761 ( .C1(n1750), .C2(n1751), .A(n1749), .B(n1752), .ZN(n1754)
         );
  NAND2_X4 U2762 ( .A1(n2281), .A2(n2280), .ZN(n2296) );
  NAND2_X4 U2763 ( .A1(net154308), .A2(net154280), .ZN(net154693) );
  NAND2_X1 U2764 ( .A1(n2773), .A2(n2772), .ZN(n2725) );
  OAI21_X4 U2765 ( .B1(n2056), .B2(n2057), .A(n1093), .ZN(n2212) );
  NOR3_X4 U2766 ( .A1(n2053), .A2(n1180), .A3(x[21]), .ZN(n2056) );
  NAND2_X4 U2767 ( .A1(n1882), .A2(n2337), .ZN(n1990) );
  NAND2_X4 U2768 ( .A1(n1920), .A2(n1919), .ZN(n1970) );
  NAND2_X4 U2769 ( .A1(n1928), .A2(n1929), .ZN(n1969) );
  NOR3_X2 U2770 ( .A1(net154802), .A2(n594), .A3(n2006), .ZN(n2007) );
  NAND2_X4 U2771 ( .A1(n2008), .A2(n2007), .ZN(n2047) );
  OAI21_X2 U2772 ( .B1(n2634), .B2(n2633), .A(n2667), .ZN(n2635) );
  NAND2_X4 U2773 ( .A1(n1536), .A2(n1537), .ZN(n1640) );
  OAI21_X4 U2774 ( .B1(n1535), .B2(n1534), .A(n1533), .ZN(n1536) );
  OAI22_X4 U2775 ( .A1(net155896), .A2(net157450), .B1(net155851), .B2(n1239), 
        .ZN(n1262) );
  INV_X8 U2776 ( .A(n1589), .ZN(n1591) );
  NAND2_X4 U2777 ( .A1(n1733), .A2(n1691), .ZN(n1881) );
  NAND2_X4 U2778 ( .A1(n1579), .A2(n1578), .ZN(n1812) );
  NAND2_X4 U2779 ( .A1(n1448), .A2(n1447), .ZN(n1545) );
  NAND2_X4 U2780 ( .A1(net155513), .A2(net157521), .ZN(n1442) );
  NAND2_X1 U2781 ( .A1(n2439), .A2(n2438), .ZN(n2440) );
  OAI21_X1 U2782 ( .B1(n1507), .B2(n628), .A(n1533), .ZN(n1508) );
  NAND2_X4 U2783 ( .A1(n1506), .A2(n1505), .ZN(n1533) );
  NAND3_X1 U2784 ( .A1(n2643), .A2(n576), .A3(n2808), .ZN(n2644) );
  NAND3_X2 U2785 ( .A1(net157542), .A2(n2130), .A3(n2085), .ZN(n2087) );
  NAND2_X4 U2786 ( .A1(n1967), .A2(n1968), .ZN(net154682) );
  NAND3_X4 U2787 ( .A1(n1980), .A2(n1979), .A3(net156073), .ZN(n1942) );
  NAND2_X4 U2788 ( .A1(net155513), .A2(net155514), .ZN(n1453) );
  INV_X32 U2789 ( .A(x[5]), .ZN(net155513) );
  NAND2_X4 U2790 ( .A1(n1624), .A2(n1637), .ZN(n1642) );
  NAND2_X1 U2791 ( .A1(n1980), .A2(n1979), .ZN(n2013) );
  NAND3_X1 U2792 ( .A1(n1709), .A2(net155665), .A3(net154943), .ZN(n1713) );
  NAND2_X4 U2793 ( .A1(net155482), .A2(net155511), .ZN(n1783) );
  INV_X32 U2794 ( .A(x[8]), .ZN(net155511) );
  INV_X8 U2795 ( .A(net154855), .ZN(net154956) );
  INV_X8 U2796 ( .A(n2818), .ZN(n2721) );
  NOR4_X4 U2797 ( .A1(n1179), .A2(n1609), .A3(n672), .A4(n1042), .ZN(n1717) );
  NAND2_X4 U2798 ( .A1(n1903), .A2(n1902), .ZN(n2341) );
  NAND2_X4 U2799 ( .A1(n2777), .A2(n2776), .ZN(n2876) );
  NAND2_X4 U2800 ( .A1(n2841), .A2(net153672), .ZN(n2752) );
  NAND4_X4 U2801 ( .A1(n2294), .A2(n2292), .A3(n2293), .A4(n2291), .ZN(n2295)
         );
  NAND2_X4 U2802 ( .A1(n1544), .A2(n1543), .ZN(n1659) );
  XNOR2_X1 U2803 ( .A(n947), .B(n1969), .ZN(n1944) );
  NAND3_X1 U2804 ( .A1(net157527), .A2(n595), .A3(net153996), .ZN(n2188) );
  NAND2_X4 U2805 ( .A1(n1431), .A2(n1496), .ZN(n1529) );
  NAND2_X4 U2806 ( .A1(y[2]), .A2(net155041), .ZN(n1559) );
  NAND3_X1 U2807 ( .A1(n883), .A2(net154481), .A3(n2187), .ZN(n2190) );
  INV_X8 U2808 ( .A(n2187), .ZN(n2314) );
  XNOR2_X1 U2809 ( .A(n1765), .B(n1891), .ZN(n1772) );
  NAND2_X1 U2810 ( .A1(net153875), .A2(n583), .ZN(n2634) );
  INV_X2 U2811 ( .A(n2408), .ZN(n2379) );
  NAND3_X2 U2812 ( .A1(n1742), .A2(n706), .A3(n1740), .ZN(n1743) );
  NAND2_X4 U2813 ( .A1(n1858), .A2(n1857), .ZN(n1863) );
  NAND2_X4 U2814 ( .A1(x[5]), .A2(n2606), .ZN(n1285) );
  NAND2_X4 U2815 ( .A1(n2582), .A2(n2581), .ZN(net153788) );
  NAND2_X4 U2816 ( .A1(n2445), .A2(n2444), .ZN(n2717) );
  NAND2_X2 U2817 ( .A1(n1965), .A2(n2345), .ZN(n2522) );
  NAND2_X4 U2818 ( .A1(n2606), .A2(x[9]), .ZN(n1572) );
  NAND2_X4 U2819 ( .A1(n2889), .A2(n2888), .ZN(n2918) );
  NAND2_X4 U2820 ( .A1(n1743), .A2(n1744), .ZN(n2514) );
  INV_X8 U2821 ( .A(n2075), .ZN(n2220) );
  NAND2_X4 U2822 ( .A1(n2074), .A2(n561), .ZN(n2075) );
  NAND2_X4 U2823 ( .A1(n2550), .A2(n2552), .ZN(n2551) );
  NAND2_X4 U2824 ( .A1(net154339), .A2(n2629), .ZN(n2549) );
  NAND2_X4 U2825 ( .A1(n2660), .A2(n2658), .ZN(n2629) );
  NAND2_X4 U2826 ( .A1(n1333), .A2(n1219), .ZN(n1587) );
  NAND2_X4 U2827 ( .A1(n1395), .A2(n1394), .ZN(n1678) );
  NAND2_X4 U2828 ( .A1(n627), .A2(n1794), .ZN(n1801) );
  NAND2_X4 U2829 ( .A1(n2555), .A2(net153986), .ZN(n2556) );
  OAI21_X2 U2830 ( .B1(n2702), .B2(n2498), .A(n2497), .ZN(n2544) );
  NAND3_X4 U2831 ( .A1(net155775), .A2(net155773), .A3(net157440), .ZN(
        net155327) );
  NAND3_X4 U2832 ( .A1(n1123), .A2(n2723), .A3(n2722), .ZN(n2769) );
  NAND2_X1 U2833 ( .A1(n1641), .A2(n1640), .ZN(n1538) );
  NAND4_X1 U2834 ( .A1(n2169), .A2(n2566), .A3(n511), .A4(n2168), .ZN(n2171)
         );
  NAND3_X2 U2835 ( .A1(n1642), .A2(n1641), .A3(n1640), .ZN(n1643) );
  NAND2_X4 U2836 ( .A1(n2429), .A2(n2395), .ZN(n2431) );
  NAND2_X4 U2837 ( .A1(n1168), .A2(n2661), .ZN(net153835) );
  NAND2_X4 U2838 ( .A1(n1967), .A2(n1968), .ZN(n2046) );
  NAND3_X4 U2839 ( .A1(n1692), .A2(n1693), .A3(n612), .ZN(n1814) );
  NAND2_X4 U2840 ( .A1(n1588), .A2(n1587), .ZN(n1693) );
  NAND2_X4 U2841 ( .A1(n2310), .A2(net157159), .ZN(n2477) );
  NAND4_X4 U2842 ( .A1(n1664), .A2(n540), .A3(n1433), .A4(n1670), .ZN(n1504)
         );
  NOR4_X4 U2843 ( .A1(x[6]), .A2(x[5]), .A3(x[8]), .A4(x[7]), .ZN(n1923) );
  OAI22_X4 U2844 ( .A1(net155885), .A2(n2052), .B1(n2112), .B2(net155855), 
        .ZN(n2084) );
  OAI21_X4 U2845 ( .B1(n1792), .B2(n1793), .A(n1941), .ZN(n1937) );
  NAND2_X4 U2846 ( .A1(n1081), .A2(n2276), .ZN(net153533) );
  XNOR2_X1 U2847 ( .A(n1960), .B(n1165), .ZN(result[18]) );
  XNOR2_X1 U2848 ( .A(n1853), .B(n806), .ZN(n1824) );
  AOI21_X1 U2849 ( .B1(n1174), .B2(net153907), .A(net156745), .ZN(
        \ddd/adder[0]/axorb ) );
  NAND2_X1 U2850 ( .A1(n1726), .A2(n978), .ZN(n1724) );
  OAI21_X1 U2851 ( .B1(n536), .B2(n1432), .A(n515), .ZN(n1460) );
  NAND2_X1 U2852 ( .A1(n1490), .A2(n515), .ZN(n1491) );
  NAND2_X1 U2853 ( .A1(n2495), .A2(n549), .ZN(n2498) );
  AOI21_X1 U2854 ( .B1(n2893), .B2(n2892), .A(n2891), .ZN(n2896) );
  NAND2_X4 U2855 ( .A1(n2525), .A2(n855), .ZN(n2720) );
  XNOR2_X1 U2856 ( .A(n2276), .B(net154339), .ZN(n2152) );
  NAND3_X2 U2857 ( .A1(n2208), .A2(n2364), .A3(net154616), .ZN(n2214) );
  NAND2_X4 U2858 ( .A1(n1604), .A2(n1062), .ZN(n1808) );
  OAI21_X2 U2859 ( .B1(net155869), .B2(n1763), .A(n1602), .ZN(n1604) );
  OAI21_X4 U2860 ( .B1(n1601), .B2(net155324), .A(n578), .ZN(n1763) );
  NOR4_X4 U2861 ( .A1(n1050), .A2(n1037), .A3(x[11]), .A4(n1554), .ZN(n1601)
         );
  NAND2_X4 U2862 ( .A1(net153930), .A2(n2589), .ZN(n2738) );
  NAND2_X4 U2863 ( .A1(n570), .A2(n1965), .ZN(n2352) );
  NAND2_X4 U2864 ( .A1(n2046), .A2(n600), .ZN(n1827) );
  NAND2_X4 U2865 ( .A1(n1813), .A2(n1812), .ZN(n1911) );
  OAI221_X4 U2866 ( .B1(net153671), .B2(n2752), .C1(n2702), .C2(n2701), .A(
        n2700), .ZN(n2703) );
  OAI211_X4 U2867 ( .C1(n1956), .C2(n1049), .A(n1955), .B(n1013), .ZN(
        net154341) );
  NAND2_X4 U2868 ( .A1(n1959), .A2(n1958), .ZN(n2289) );
  NAND2_X4 U2869 ( .A1(n935), .A2(n2750), .ZN(net153669) );
  AOI211_X4 U2870 ( .C1(n2721), .C2(n1029), .A(net153881), .B(n2628), .ZN(
        n2641) );
  NAND2_X4 U2871 ( .A1(n2626), .A2(n2625), .ZN(n2809) );
  NAND3_X1 U2872 ( .A1(n841), .A2(n2159), .A3(n805), .ZN(n2155) );
  INV_X8 U2873 ( .A(net154578), .ZN(net154031) );
  NAND2_X1 U2874 ( .A1(n2437), .A2(n686), .ZN(n2439) );
  NAND2_X1 U2875 ( .A1(n2065), .A2(net154038), .ZN(n2040) );
  INV_X32 U2876 ( .A(y[1]), .ZN(net155041) );
  NAND2_X4 U2877 ( .A1(y[0]), .A2(net155041), .ZN(n2533) );
  NAND2_X4 U2878 ( .A1(y[1]), .A2(net155739), .ZN(net153818) );
  NAND2_X4 U2879 ( .A1(n2508), .A2(net154055), .ZN(net153828) );
  NAND3_X4 U2880 ( .A1(y[0]), .A2(net155041), .A3(x[1]), .ZN(n1188) );
  NAND2_X2 U2881 ( .A1(net155777), .A2(net155819), .ZN(n1187) );
  NAND2_X2 U2882 ( .A1(n1188), .A2(n1187), .ZN(n1185) );
  INV_X4 U2883 ( .A(n1559), .ZN(n1196) );
  INV_X4 U2884 ( .A(n1184), .ZN(n1915) );
  NAND3_X4 U2885 ( .A1(y[1]), .A2(net155739), .A3(x[1]), .ZN(net155799) );
  OAI21_X4 U2886 ( .B1(x[1]), .B2(x[0]), .A(x[2]), .ZN(n1213) );
  NAND3_X4 U2887 ( .A1(y[0]), .A2(net155041), .A3(x[2]), .ZN(n1199) );
  XNOR2_X2 U2888 ( .A(net155815), .B(n1186), .ZN(n1192) );
  INV_X4 U2889 ( .A(n1187), .ZN(n1191) );
  INV_X4 U2890 ( .A(n1188), .ZN(n1190) );
  OAI21_X4 U2891 ( .B1(n1191), .B2(n1190), .A(n713), .ZN(n1220) );
  NAND2_X2 U2892 ( .A1(n1193), .A2(n1223), .ZN(n1227) );
  NAND2_X2 U2893 ( .A1(n1194), .A2(n1227), .ZN(n1195) );
  INV_X4 U2894 ( .A(n1195), .ZN(n1205) );
  OAI21_X4 U2895 ( .B1(net155847), .B2(net153769), .A(net157416), .ZN(n1204)
         );
  XNOR2_X2 U2896 ( .A(n1205), .B(n1204), .ZN(result[2]) );
  OAI21_X4 U2897 ( .B1(x[1]), .B2(x[0]), .A(x[2]), .ZN(n1197) );
  NOR2_X4 U2898 ( .A1(x[3]), .A2(x[0]), .ZN(n1209) );
  OAI21_X4 U2899 ( .B1(n1223), .B2(n1201), .A(n1245), .ZN(n1202) );
  XNOR2_X2 U2900 ( .A(n1203), .B(n1202), .ZN(n1233) );
  INV_X4 U2901 ( .A(n1204), .ZN(n1206) );
  INV_X4 U2902 ( .A(n1237), .ZN(n1208) );
  INV_X4 U2903 ( .A(y[4]), .ZN(net155791) );
  INV_X4 U2904 ( .A(n1207), .ZN(n1238) );
  XNOR2_X2 U2905 ( .A(n1208), .B(n1238), .ZN(result[3]) );
  INV_X4 U2906 ( .A(net155732), .ZN(net155780) );
  INV_X4 U2907 ( .A(net155697), .ZN(net155781) );
  OAI21_X4 U2908 ( .B1(net155780), .B2(net155781), .A(net155782), .ZN(n1255)
         );
  NAND2_X2 U2909 ( .A1(n1217), .A2(n1216), .ZN(n1218) );
  NAND2_X2 U2910 ( .A1(n1228), .A2(n1288), .ZN(n1257) );
  NAND2_X2 U2911 ( .A1(n1227), .A2(n1226), .ZN(n1229) );
  XNOR2_X2 U2912 ( .A(n1229), .B(n598), .ZN(n1231) );
  NAND2_X2 U2913 ( .A1(n1265), .A2(n1264), .ZN(n1274) );
  INV_X4 U2914 ( .A(n1274), .ZN(n1235) );
  XNOR2_X2 U2915 ( .A(n1236), .B(n1235), .ZN(n1270) );
  NAND2_X2 U2916 ( .A1(n1238), .A2(n1237), .ZN(n1269) );
  OAI22_X2 U2917 ( .A1(n2705), .A2(net157451), .B1(net155827), .B2(n1239), 
        .ZN(n1316) );
  NOR3_X4 U2918 ( .A1(x[0]), .A2(x[2]), .A3(x[1]), .ZN(n1240) );
  NAND2_X2 U2919 ( .A1(x[4]), .A2(net155884), .ZN(n1242) );
  XNOR2_X2 U2920 ( .A(n1310), .B(net155657), .ZN(n1254) );
  NAND2_X2 U2921 ( .A1(n1246), .A2(n1288), .ZN(n1308) );
  INV_X4 U2922 ( .A(n1308), .ZN(n1248) );
  NAND2_X2 U2923 ( .A1(n1248), .A2(n557), .ZN(n1252) );
  NAND2_X2 U2924 ( .A1(n1250), .A2(n1249), .ZN(n1251) );
  INV_X4 U2925 ( .A(n1309), .ZN(n1261) );
  INV_X4 U2926 ( .A(n1257), .ZN(n1259) );
  XNOR2_X2 U2927 ( .A(n1261), .B(n1260), .ZN(n1263) );
  NAND2_X2 U2928 ( .A1(n1263), .A2(n1262), .ZN(n1345) );
  INV_X4 U2929 ( .A(n1265), .ZN(n1266) );
  OAI21_X4 U2930 ( .B1(n1267), .B2(n1266), .A(n923), .ZN(n1344) );
  XNOR2_X2 U2931 ( .A(n1268), .B(n1315), .ZN(n1320) );
  INV_X4 U2932 ( .A(n1269), .ZN(n1271) );
  INV_X4 U2933 ( .A(n1272), .ZN(n1314) );
  XNOR2_X2 U2934 ( .A(n1278), .B(n1277), .ZN(result[5]) );
  NAND3_X4 U2935 ( .A1(n1291), .A2(n510), .A3(n1412), .ZN(n1471) );
  NAND2_X2 U2936 ( .A1(n1471), .A2(n1293), .ZN(n1340) );
  INV_X4 U2937 ( .A(n1294), .ZN(n1295) );
  NOR2_X4 U2938 ( .A1(n1295), .A2(net155592), .ZN(n1302) );
  NOR2_X4 U2939 ( .A1(x[6]), .A2(x[5]), .ZN(n1297) );
  NOR2_X4 U2940 ( .A1(x[4]), .A2(x[3]), .ZN(n1296) );
  NAND2_X2 U2941 ( .A1(x[6]), .A2(n2606), .ZN(n1300) );
  OAI21_X4 U2942 ( .B1(n1302), .B2(n1301), .A(n1300), .ZN(n1407) );
  XNOR2_X2 U2943 ( .A(n1332), .B(n1331), .ZN(n1339) );
  OAI22_X2 U2944 ( .A1(net155896), .A2(net155645), .B1(net155839), .B2(n1321), 
        .ZN(n1341) );
  XNOR2_X2 U2945 ( .A(n1339), .B(n1341), .ZN(n1305) );
  XNOR2_X2 U2946 ( .A(n1340), .B(n1305), .ZN(n1350) );
  XNOR2_X2 U2947 ( .A(n1352), .B(n1350), .ZN(n1313) );
  NAND2_X2 U2948 ( .A1(n1312), .A2(net155657), .ZN(n1360) );
  NAND2_X2 U2949 ( .A1(n1361), .A2(n1360), .ZN(n1351) );
  XNOR2_X2 U2950 ( .A(n1313), .B(n1351), .ZN(n1517) );
  NOR2_X4 U2951 ( .A1(n1314), .A2(n532), .ZN(n1319) );
  NAND2_X2 U2952 ( .A1(n1317), .A2(n1316), .ZN(n1318) );
  OAI21_X4 U2953 ( .B1(n1320), .B2(n1319), .A(n1318), .ZN(n1349) );
  OAI22_X2 U2954 ( .A1(n2705), .A2(net155665), .B1(net155827), .B2(n1321), 
        .ZN(n1356) );
  NAND2_X2 U2955 ( .A1(x[6]), .A2(net155884), .ZN(n1323) );
  NOR2_X4 U2956 ( .A1(n1324), .A2(n1116), .ZN(n1325) );
  INV_X4 U2957 ( .A(n1328), .ZN(n1330) );
  OAI21_X4 U2958 ( .B1(n1330), .B2(n1329), .A(n1407), .ZN(n1403) );
  INV_X4 U2959 ( .A(x[5]), .ZN(net155624) );
  INV_X4 U2960 ( .A(n1360), .ZN(n1347) );
  AOI21_X4 U2961 ( .B1(n1344), .B2(n1345), .A(n1343), .ZN(n1346) );
  XNOR2_X2 U2962 ( .A(n1348), .B(n1355), .ZN(n1519) );
  XNOR2_X2 U2963 ( .A(n1351), .B(n603), .ZN(n1353) );
  XNOR2_X2 U2964 ( .A(n1358), .B(n1354), .ZN(result[7]) );
  INV_X4 U2965 ( .A(n1354), .ZN(n1359) );
  OAI21_X4 U2966 ( .B1(n1359), .B2(n1358), .A(n1523), .ZN(n1392) );
  INV_X4 U2967 ( .A(n1392), .ZN(n1388) );
  INV_X4 U2968 ( .A(n1493), .ZN(n1362) );
  AOI21_X4 U2969 ( .B1(n1364), .B2(n1363), .A(n1362), .ZN(n1368) );
  OAI21_X4 U2970 ( .B1(n1368), .B2(n1396), .A(n1494), .ZN(n1526) );
  INV_X4 U2971 ( .A(x[6]), .ZN(net155592) );
  NAND2_X2 U2972 ( .A1(x[8]), .A2(n2606), .ZN(n1375) );
  INV_X4 U2973 ( .A(n1471), .ZN(n1379) );
  OAI21_X4 U2974 ( .B1(n1326), .B2(net155869), .A(n1382), .ZN(n1402) );
  XNOR2_X2 U2975 ( .A(n1385), .B(n1141), .ZN(n1525) );
  INV_X4 U2976 ( .A(n1389), .ZN(n1387) );
  NAND2_X2 U2977 ( .A1(x[5]), .A2(n1183), .ZN(n1386) );
  FA_X1 U2978 ( .A(n1388), .B(n1387), .CI(n1527), .S(result[8]) );
  NAND2_X2 U2979 ( .A1(n1389), .A2(n1527), .ZN(n1490) );
  XNOR2_X2 U2980 ( .A(n1390), .B(n1526), .ZN(n1522) );
  NAND2_X2 U2981 ( .A1(n1392), .A2(n1391), .ZN(n1489) );
  NAND3_X4 U2982 ( .A1(n1494), .A2(n539), .A3(n1396), .ZN(n1433) );
  NAND3_X2 U2983 ( .A1(n540), .A2(n1670), .A3(n1433), .ZN(n1430) );
  INV_X4 U2984 ( .A(n1398), .ZN(n1400) );
  OAI21_X4 U2985 ( .B1(n1401), .B2(n1400), .A(n1399), .ZN(n1571) );
  NAND2_X2 U2986 ( .A1(x[8]), .A2(net155884), .ZN(n1416) );
  INV_X4 U2987 ( .A(n1574), .ZN(n1419) );
  AOI21_X4 U2988 ( .B1(n1596), .B2(n842), .A(n1419), .ZN(n1420) );
  XNOR2_X2 U2989 ( .A(n1577), .B(n1420), .ZN(n1422) );
  NAND3_X2 U2990 ( .A1(n575), .A2(n992), .A3(n934), .ZN(n1424) );
  XNOR2_X2 U2991 ( .A(n1434), .B(n1435), .ZN(n1497) );
  NAND2_X2 U2992 ( .A1(x[6]), .A2(n1183), .ZN(n1426) );
  XNOR2_X2 U2993 ( .A(n1428), .B(n1496), .ZN(n1432) );
  INV_X4 U2994 ( .A(n1432), .ZN(n1429) );
  XNOR2_X2 U2995 ( .A(n536), .B(n1429), .ZN(result[9]) );
  XNOR2_X2 U2996 ( .A(n1430), .B(n1497), .ZN(n1431) );
  XNOR2_X2 U2997 ( .A(n1434), .B(n1435), .ZN(n1664) );
  OAI21_X4 U2998 ( .B1(n1596), .B2(net155869), .A(n842), .ZN(n1438) );
  OAI21_X4 U2999 ( .B1(n1441), .B2(n1440), .A(n1439), .ZN(n1463) );
  NOR2_X4 U3000 ( .A1(x[10]), .A2(x[9]), .ZN(n1608) );
  NOR2_X4 U3001 ( .A1(x[6]), .A2(x[5]), .ZN(n1548) );
  NAND2_X2 U3002 ( .A1(n1449), .A2(n1545), .ZN(n1450) );
  NAND2_X2 U3003 ( .A1(x[10]), .A2(n2606), .ZN(n1466) );
  NAND3_X2 U3004 ( .A1(n1450), .A2(n1467), .A3(n1466), .ZN(n1452) );
  NAND2_X2 U3005 ( .A1(n1466), .A2(net155873), .ZN(n1451) );
  NOR2_X4 U3006 ( .A1(x[1]), .A2(x[0]), .ZN(n1455) );
  NOR3_X4 U3007 ( .A1(x[2]), .A2(x[4]), .A3(x[3]), .ZN(n1454) );
  INV_X4 U3008 ( .A(x[8]), .ZN(net155484) );
  INV_X4 U3009 ( .A(n1464), .ZN(n1656) );
  XNOR2_X2 U3010 ( .A(n1463), .B(n1665), .ZN(n1617) );
  XNOR2_X2 U3011 ( .A(n1459), .B(n1458), .ZN(n1500) );
  INV_X4 U3012 ( .A(n1510), .ZN(n1513) );
  NAND2_X2 U3013 ( .A1(n1539), .A2(n1541), .ZN(n1512) );
  AOI21_X2 U3014 ( .B1(n1588), .B2(n1471), .A(n921), .ZN(n1476) );
  NAND3_X2 U3015 ( .A1(n1476), .A2(n1474), .A3(n1475), .ZN(n1477) );
  NAND2_X2 U3016 ( .A1(x[10]), .A2(net155884), .ZN(n1481) );
  NOR2_X4 U3017 ( .A1(n543), .A2(net155857), .ZN(n1479) );
  INV_X4 U3018 ( .A(n1695), .ZN(n1700) );
  NAND2_X2 U3019 ( .A1(x[11]), .A2(n2606), .ZN(n1568) );
  INV_X4 U3020 ( .A(n1568), .ZN(n1486) );
  XNOR2_X2 U3021 ( .A(n1484), .B(x[11]), .ZN(n1567) );
  NAND2_X2 U3022 ( .A1(n1568), .A2(net155873), .ZN(n1485) );
  INV_X4 U3023 ( .A(n1699), .ZN(n1487) );
  XNOR2_X2 U3024 ( .A(n1700), .B(n1487), .ZN(n1590) );
  INV_X4 U3025 ( .A(x[9]), .ZN(net155446) );
  OAI22_X2 U3026 ( .A1(net155896), .A2(net155446), .B1(n1596), .B2(net155841), 
        .ZN(n1543) );
  XNOR2_X2 U3027 ( .A(n1590), .B(n1543), .ZN(n1488) );
  XNOR2_X2 U3028 ( .A(n1542), .B(n1488), .ZN(n1540) );
  INV_X4 U3029 ( .A(n1489), .ZN(n1492) );
  NAND2_X2 U3030 ( .A1(n1494), .A2(n1493), .ZN(n1675) );
  INV_X4 U3031 ( .A(n1494), .ZN(n1677) );
  XNOR2_X2 U3032 ( .A(n1499), .B(n1498), .ZN(n1503) );
  INV_X4 U3033 ( .A(n1500), .ZN(n1501) );
  OAI21_X4 U3034 ( .B1(n1503), .B2(n1502), .A(n1501), .ZN(n1534) );
  FA_X1 U3035 ( .A(n1513), .B(n1509), .CI(n1508), .S(result[11]) );
  NAND2_X2 U3036 ( .A1(n1511), .A2(n1510), .ZN(n1641) );
  XNOR2_X2 U3037 ( .A(n1619), .B(n1513), .ZN(n1514) );
  XNOR2_X2 U3038 ( .A(n1515), .B(n1514), .ZN(n1537) );
  INV_X4 U3039 ( .A(n1516), .ZN(n1521) );
  OAI21_X4 U3040 ( .B1(n1520), .B2(n1521), .A(n1519), .ZN(n1524) );
  NOR2_X4 U3041 ( .A1(n1532), .A2(n1531), .ZN(n1535) );
  INV_X4 U3042 ( .A(n1538), .ZN(n1626) );
  XOR2_X2 U3043 ( .A(n1542), .B(n555), .Z(n1544) );
  NAND2_X2 U3044 ( .A1(x[10]), .A2(net153769), .ZN(n1547) );
  OAI21_X4 U3045 ( .B1(net155839), .B2(n1613), .A(n1547), .ZN(n1647) );
  NOR2_X4 U3046 ( .A1(x[10]), .A2(x[9]), .ZN(n1549) );
  NOR2_X4 U3047 ( .A1(x[11]), .A2(x[4]), .ZN(n1551) );
  NOR2_X4 U3048 ( .A1(x[12]), .A2(x[3]), .ZN(n1550) );
  NOR2_X4 U3049 ( .A1(x[8]), .A2(x[7]), .ZN(n1552) );
  INV_X4 U3050 ( .A(n1552), .ZN(n1597) );
  NOR2_X4 U3051 ( .A1(x[10]), .A2(x[9]), .ZN(n1787) );
  NAND3_X4 U3052 ( .A1(y[0]), .A2(net155041), .A3(x[12]), .ZN(n1602) );
  NAND2_X2 U3053 ( .A1(x[12]), .A2(n1602), .ZN(n1556) );
  NAND2_X2 U3054 ( .A1(n1602), .A2(net155873), .ZN(n1555) );
  NOR2_X4 U3055 ( .A1(n1558), .A2(n1557), .ZN(n1694) );
  NAND2_X2 U3056 ( .A1(x[11]), .A2(net155884), .ZN(n1565) );
  NOR3_X4 U3057 ( .A1(net155367), .A2(n1561), .A3(n1560), .ZN(n1562) );
  XNOR2_X2 U3058 ( .A(n1562), .B(n1563), .ZN(n1564) );
  XNOR2_X2 U3059 ( .A(n1694), .B(n1566), .ZN(n1701) );
  OAI21_X4 U3060 ( .B1(n1723), .B2(net155869), .A(n1568), .ZN(n1696) );
  INV_X4 U3061 ( .A(n1572), .ZN(n1573) );
  INV_X4 U3062 ( .A(n1583), .ZN(n1584) );
  NAND3_X4 U3063 ( .A1(n1693), .A2(n1692), .A3(n612), .ZN(n1589) );
  OAI21_X4 U3064 ( .B1(n1592), .B2(n1591), .A(n555), .ZN(n1618) );
  XNOR2_X2 U3065 ( .A(n1594), .B(n680), .ZN(n1623) );
  NAND2_X2 U3066 ( .A1(x[9]), .A2(n1183), .ZN(n1595) );
  XNOR2_X2 U3067 ( .A(n1626), .B(n1622), .ZN(result[12]) );
  INV_X4 U3068 ( .A(n1618), .ZN(n1686) );
  INV_X4 U3069 ( .A(x[12]), .ZN(net155324) );
  NOR2_X4 U3070 ( .A1(n1609), .A2(n1597), .ZN(n1600) );
  NAND2_X2 U3071 ( .A1(n1684), .A2(n857), .ZN(n1606) );
  NAND2_X2 U3072 ( .A1(n1687), .A2(n857), .ZN(n1605) );
  OAI21_X4 U3073 ( .B1(n1606), .B2(n1686), .A(n1605), .ZN(n1612) );
  NAND2_X2 U3074 ( .A1(x[12]), .A2(net155884), .ZN(n1607) );
  XNOR2_X2 U3075 ( .A(n1717), .B(x[13]), .ZN(n1759) );
  INV_X4 U3076 ( .A(x[11]), .ZN(net155310) );
  OAI22_X2 U3077 ( .A1(net155896), .A2(net155310), .B1(n829), .B2(net155841), 
        .ZN(n1691) );
  INV_X4 U3078 ( .A(n1691), .ZN(n1735) );
  INV_X4 U3079 ( .A(x[10]), .ZN(n1614) );
  OAI22_X2 U3080 ( .A1(n2705), .A2(n1614), .B1(net155827), .B2(n1613), .ZN(
        n1634) );
  INV_X4 U3081 ( .A(n1634), .ZN(n1615) );
  XNOR2_X2 U3082 ( .A(n1616), .B(n1615), .ZN(n1639) );
  NAND2_X2 U3083 ( .A1(n1648), .A2(n1647), .ZN(n1653) );
  NAND3_X2 U3084 ( .A1(n1630), .A2(n1086), .A3(n534), .ZN(n1621) );
  NAND2_X2 U3085 ( .A1(n1629), .A2(n1086), .ZN(n1620) );
  XNOR2_X2 U3086 ( .A(n1639), .B(n1638), .ZN(n1628) );
  INV_X4 U3087 ( .A(n1622), .ZN(n1625) );
  INV_X4 U3088 ( .A(n1623), .ZN(n1624) );
  XNOR2_X2 U3089 ( .A(n1628), .B(n1627), .ZN(result[13]) );
  INV_X4 U3090 ( .A(n1629), .ZN(n1632) );
  NAND2_X2 U3091 ( .A1(n534), .A2(n1630), .ZN(n1631) );
  INV_X4 U3092 ( .A(n1653), .ZN(n1738) );
  AOI21_X4 U3093 ( .B1(n1632), .B2(n1631), .A(n1738), .ZN(n1633) );
  NAND2_X2 U3094 ( .A1(n1635), .A2(n1634), .ZN(n1726) );
  FA_X1 U3095 ( .A(n1637), .B(n680), .CI(n1594), .S(n1645) );
  OAI21_X4 U3096 ( .B1(n1650), .B2(n1079), .A(n1649), .ZN(n1651) );
  INV_X4 U3097 ( .A(n1652), .ZN(n1654) );
  XNOR2_X2 U3098 ( .A(n1656), .B(n1655), .ZN(n1658) );
  OAI21_X4 U3099 ( .B1(n1661), .B2(n1660), .A(n1659), .ZN(n1662) );
  NAND3_X4 U3100 ( .A1(n1741), .A2(n1663), .A3(n1736), .ZN(n1767) );
  INV_X4 U3101 ( .A(n1664), .ZN(n1673) );
  INV_X4 U3102 ( .A(n1670), .ZN(n1671) );
  NOR3_X4 U3103 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1769) );
  NOR2_X4 U3104 ( .A1(n1676), .A2(n1675), .ZN(n1680) );
  OAI21_X4 U3105 ( .B1(n1680), .B2(n1679), .A(n539), .ZN(n1768) );
  INV_X4 U3106 ( .A(n1684), .ZN(n1685) );
  NOR2_X4 U3107 ( .A1(n1686), .A2(n1685), .ZN(n1688) );
  OAI21_X4 U3108 ( .B1(n1688), .B2(n1687), .A(n857), .ZN(n1690) );
  NAND2_X2 U3109 ( .A1(n538), .A2(n1881), .ZN(n1721) );
  NAND3_X2 U3110 ( .A1(n1695), .A2(n1694), .A3(n1696), .ZN(n1809) );
  NOR2_X2 U3111 ( .A1(n856), .A2(n1697), .ZN(n1698) );
  NAND2_X2 U3112 ( .A1(n1698), .A2(n1812), .ZN(n1750) );
  NAND2_X2 U3113 ( .A1(n1700), .A2(n1699), .ZN(n1702) );
  NAND2_X2 U3114 ( .A1(n1147), .A2(n1830), .ZN(n1703) );
  INV_X4 U3115 ( .A(n1705), .ZN(n1706) );
  OAI21_X4 U3116 ( .B1(n1707), .B2(n1706), .A(n711), .ZN(n1886) );
  NOR2_X4 U3117 ( .A1(x[13]), .A2(x[11]), .ZN(n1709) );
  NOR2_X4 U3118 ( .A1(x[12]), .A2(x[3]), .ZN(n1781) );
  OAI21_X4 U3119 ( .B1(n1713), .B2(n1712), .A(x[14]), .ZN(n1755) );
  XNOR2_X2 U3120 ( .A(n1717), .B(x[13]), .ZN(n1718) );
  XNOR2_X2 U3121 ( .A(n930), .B(n1794), .ZN(n1748) );
  INV_X4 U3122 ( .A(n1728), .ZN(n1719) );
  XNOR2_X2 U3123 ( .A(n1889), .B(n1719), .ZN(n1720) );
  XNOR2_X2 U3124 ( .A(n1721), .B(n898), .ZN(n1865) );
  NAND2_X2 U3125 ( .A1(x[11]), .A2(n1183), .ZN(n1722) );
  INV_X4 U3126 ( .A(n1726), .ZN(n1870) );
  XNOR2_X2 U3127 ( .A(n1890), .B(n831), .ZN(n1729) );
  NAND2_X2 U3128 ( .A1(n1731), .A2(n1730), .ZN(n1732) );
  AOI21_X2 U3129 ( .B1(n1732), .B2(n1881), .A(n898), .ZN(n1744) );
  INV_X4 U3130 ( .A(n1810), .ZN(n1888) );
  NAND2_X2 U3131 ( .A1(net155884), .A2(x[14]), .ZN(n1756) );
  OAI21_X4 U3132 ( .B1(net155855), .B2(n1847), .A(n1756), .ZN(n1798) );
  NAND2_X2 U3133 ( .A1(x[15]), .A2(n2606), .ZN(n1757) );
  OAI21_X4 U3134 ( .B1(n958), .B2(net155869), .A(n1757), .ZN(n1797) );
  XNOR2_X2 U3135 ( .A(n1798), .B(n1797), .ZN(n1835) );
  NAND2_X2 U3136 ( .A1(x[13]), .A2(net153769), .ZN(n1760) );
  XNOR2_X2 U3137 ( .A(n1761), .B(n803), .ZN(n1856) );
  NAND2_X2 U3138 ( .A1(x[12]), .A2(n1183), .ZN(n1762) );
  XNOR2_X2 U3139 ( .A(n1764), .B(n2024), .ZN(result[15]) );
  INV_X4 U3140 ( .A(n1766), .ZN(n1828) );
  NOR2_X4 U3141 ( .A1(n1771), .A2(n1770), .ZN(n1956) );
  NAND2_X2 U3142 ( .A1(x[14]), .A2(net153769), .ZN(n1775) );
  XNOR2_X2 U3143 ( .A(x[15]), .B(n1776), .ZN(n1778) );
  NAND2_X2 U3144 ( .A1(x[15]), .A2(net155884), .ZN(n1777) );
  OAI21_X4 U3145 ( .B1(n1778), .B2(net155857), .A(n1777), .ZN(n1837) );
  INV_X4 U3146 ( .A(x[16]), .ZN(n1793) );
  INV_X4 U3147 ( .A(x[11]), .ZN(net155112) );
  INV_X4 U3148 ( .A(n1784), .ZN(n1785) );
  NOR2_X4 U3149 ( .A1(x[12]), .A2(x[11]), .ZN(n1788) );
  INV_X4 U3150 ( .A(n1798), .ZN(n1799) );
  OAI21_X4 U3151 ( .B1(n1888), .B2(n1831), .A(n1803), .ZN(n1806) );
  NAND3_X2 U3152 ( .A1(n1830), .A2(n1804), .A3(n1803), .ZN(n1805) );
  NOR2_X4 U3153 ( .A1(n942), .A2(n1811), .ZN(n1813) );
  INV_X4 U3154 ( .A(x[13]), .ZN(n1818) );
  INV_X4 U3155 ( .A(n1823), .ZN(n1819) );
  INV_X4 U3156 ( .A(n2028), .ZN(n1822) );
  INV_X4 U3157 ( .A(n1821), .ZN(n1825) );
  XNOR2_X2 U3158 ( .A(n1822), .B(n1825), .ZN(result[16]) );
  OAI21_X4 U3159 ( .B1(n1874), .B2(n1873), .A(n1872), .ZN(n2256) );
  INV_X4 U3160 ( .A(n562), .ZN(n1834) );
  INV_X4 U3161 ( .A(x[15]), .ZN(n1839) );
  NAND3_X4 U3162 ( .A1(y[0]), .A2(net155041), .A3(x[17]), .ZN(n1904) );
  NAND2_X2 U3163 ( .A1(x[17]), .A2(n1904), .ZN(n1842) );
  XNOR2_X2 U3164 ( .A(n1843), .B(n1842), .ZN(n1972) );
  NAND2_X2 U3165 ( .A1(n1904), .A2(net155873), .ZN(n1973) );
  NAND2_X2 U3166 ( .A1(x[16]), .A2(net155884), .ZN(n1844) );
  OAI21_X4 U3167 ( .B1(net155855), .B2(n1937), .A(n1844), .ZN(n1971) );
  XNOR2_X2 U3168 ( .A(n1971), .B(n1845), .ZN(net154968) );
  XNOR2_X2 U3169 ( .A(n1901), .B(n1846), .ZN(n1994) );
  INV_X4 U3170 ( .A(x[14]), .ZN(n1848) );
  INV_X4 U3171 ( .A(n1876), .ZN(n1849) );
  XNOR2_X2 U3172 ( .A(n1850), .B(n1849), .ZN(n2255) );
  XNOR2_X2 U3173 ( .A(n1875), .B(n2255), .ZN(n2034) );
  XNOR2_X2 U3174 ( .A(n1851), .B(n2034), .ZN(result[17]) );
  INV_X4 U3175 ( .A(n2034), .ZN(n2169) );
  XNOR2_X2 U3176 ( .A(n1853), .B(n1852), .ZN(n1867) );
  INV_X4 U3177 ( .A(n1867), .ZN(n1859) );
  INV_X4 U3178 ( .A(n1854), .ZN(n1860) );
  INV_X4 U3179 ( .A(n1855), .ZN(n1858) );
  NAND3_X2 U3180 ( .A1(n1860), .A2(n1859), .A3(n1863), .ZN(n1861) );
  NAND3_X2 U3181 ( .A1(n1861), .A2(n2026), .A3(n1862), .ZN(n2265) );
  INV_X4 U3182 ( .A(n1863), .ZN(n1868) );
  OAI21_X4 U3183 ( .B1(n1871), .B2(n1870), .A(n1869), .ZN(n2761) );
  XNOR2_X2 U3184 ( .A(n2256), .B(n1013), .ZN(n1877) );
  NAND4_X2 U3185 ( .A1(n1881), .A2(n1125), .A3(n1882), .A4(n2337), .ZN(n2219)
         );
  INV_X4 U3186 ( .A(n1885), .ZN(n1989) );
  NOR3_X4 U3187 ( .A1(n1990), .A2(n2342), .A3(n1989), .ZN(n1899) );
  INV_X4 U3188 ( .A(n1891), .ZN(n1892) );
  XNOR2_X2 U3189 ( .A(n1146), .B(n1892), .ZN(n1893) );
  XNOR2_X2 U3190 ( .A(n1894), .B(n1893), .ZN(n1896) );
  NOR3_X4 U3191 ( .A1(n1996), .A2(n2340), .A3(n1952), .ZN(n1898) );
  OAI211_X2 U3192 ( .C1(n1956), .C2(n1049), .A(n1900), .B(n1013), .ZN(n1936)
         );
  NAND2_X2 U3193 ( .A1(n1936), .A2(n1027), .ZN(n1933) );
  OAI21_X4 U3194 ( .B1(n572), .B2(net155869), .A(n1904), .ZN(n1905) );
  INV_X4 U3195 ( .A(net154877), .ZN(net154964) );
  NOR2_X4 U3196 ( .A1(net154964), .A2(n1910), .ZN(n1909) );
  XNOR2_X2 U3197 ( .A(n1917), .B(n1918), .ZN(n1920) );
  NAND2_X2 U3198 ( .A1(n1947), .A2(net155855), .ZN(n1919) );
  NOR2_X4 U3199 ( .A1(x[16]), .A2(x[15]), .ZN(n1922) );
  NOR2_X4 U3200 ( .A1(x[10]), .A2(x[9]), .ZN(n1921) );
  AOI21_X4 U3201 ( .B1(n2012), .B2(n1925), .A(n1924), .ZN(n1929) );
  NOR2_X4 U3202 ( .A1(x[17]), .A2(net155869), .ZN(n1927) );
  INV_X4 U3203 ( .A(n1944), .ZN(n1935) );
  NAND2_X2 U3204 ( .A1(x[16]), .A2(net153769), .ZN(n1930) );
  XNOR2_X2 U3205 ( .A(n1935), .B(n2335), .ZN(n1931) );
  NAND2_X2 U3206 ( .A1(x[15]), .A2(n1183), .ZN(n1932) );
  INV_X4 U3207 ( .A(n2282), .ZN(n2257) );
  XNOR2_X2 U3208 ( .A(n1933), .B(n1965), .ZN(n2283) );
  NAND2_X2 U3209 ( .A1(n969), .A2(n1936), .ZN(n1964) );
  NAND2_X2 U3210 ( .A1(n1964), .A2(n1089), .ZN(n1950) );
  NAND2_X2 U3211 ( .A1(x[17]), .A2(net153769), .ZN(n1938) );
  NAND2_X2 U3212 ( .A1(x[19]), .A2(n2606), .ZN(net154880) );
  NAND2_X2 U3213 ( .A1(x[18]), .A2(net155884), .ZN(n1943) );
  NAND2_X2 U3214 ( .A1(x[17]), .A2(x[18]), .ZN(n1939) );
  NAND3_X2 U3215 ( .A1(n1946), .A2(n1945), .A3(n1043), .ZN(n2353) );
  NOR3_X4 U3216 ( .A1(n1996), .A2(n2340), .A3(n1952), .ZN(n1953) );
  NAND2_X2 U3217 ( .A1(n2016), .A2(n1089), .ZN(n1957) );
  XNOR2_X2 U3218 ( .A(n1957), .B(net157139), .ZN(n1959) );
  INV_X4 U3219 ( .A(n1964), .ZN(n1966) );
  OAI21_X4 U3220 ( .B1(n1975), .B2(n1974), .A(net154285), .ZN(net154815) );
  INV_X4 U3221 ( .A(net154867), .ZN(net154827) );
  NAND2_X2 U3222 ( .A1(net154827), .A2(net154826), .ZN(n1976) );
  INV_X4 U3223 ( .A(x[19]), .ZN(net154863) );
  INV_X4 U3224 ( .A(x[20]), .ZN(net154852) );
  INV_X4 U3225 ( .A(x[12]), .ZN(net154861) );
  NAND2_X2 U3226 ( .A1(x[18]), .A2(net153769), .ZN(n1981) );
  OAI21_X4 U3227 ( .B1(net155839), .B2(n2013), .A(n1981), .ZN(net154534) );
  INV_X4 U3228 ( .A(net154534), .ZN(net154848) );
  XNOR2_X2 U3229 ( .A(n1999), .B(n1998), .ZN(n2154) );
  INV_X4 U3230 ( .A(n2154), .ZN(n2066) );
  NAND2_X2 U3231 ( .A1(x[17]), .A2(n1183), .ZN(n1982) );
  INV_X4 U3232 ( .A(n2270), .ZN(n1983) );
  XNOR2_X2 U3233 ( .A(n2066), .B(n1983), .ZN(n2286) );
  NAND2_X2 U3234 ( .A1(n2285), .A2(n2284), .ZN(net154842) );
  NOR2_X4 U3235 ( .A1(net154829), .A2(net154828), .ZN(n1997) );
  OAI21_X4 U3236 ( .B1(n1997), .B2(net154826), .A(net154827), .ZN(net154824)
         );
  XNOR2_X2 U3237 ( .A(n1999), .B(n1998), .ZN(net154028) );
  NAND2_X2 U3238 ( .A1(n2065), .A2(n561), .ZN(n2017) );
  INV_X4 U3239 ( .A(n2003), .ZN(n2085) );
  XNOR2_X2 U3240 ( .A(x[21]), .B(n2047), .ZN(n2011) );
  NAND2_X2 U3241 ( .A1(x[21]), .A2(n2606), .ZN(n2049) );
  INV_X4 U3242 ( .A(n2049), .ZN(n2009) );
  NOR2_X4 U3243 ( .A1(n692), .A2(n2009), .ZN(n2010) );
  INV_X4 U3244 ( .A(net154788), .ZN(net154719) );
  INV_X4 U3245 ( .A(x[18]), .ZN(net154784) );
  INV_X4 U3246 ( .A(n2022), .ZN(n2277) );
  INV_X4 U3247 ( .A(n2016), .ZN(n2070) );
  NAND2_X2 U3248 ( .A1(n2134), .A2(n2018), .ZN(n2020) );
  NAND2_X2 U3249 ( .A1(n2018), .A2(n2017), .ZN(n2019) );
  XNOR2_X2 U3250 ( .A(net154606), .B(net154533), .ZN(n2080) );
  XNOR2_X2 U3251 ( .A(n2021), .B(n2080), .ZN(n2278) );
  INV_X4 U3252 ( .A(n2278), .ZN(n2023) );
  INV_X4 U3253 ( .A(n2170), .ZN(n2178) );
  INV_X4 U3254 ( .A(n1764), .ZN(n2025) );
  NOR3_X4 U3255 ( .A1(n2025), .A2(n2024), .A3(n2028), .ZN(n2030) );
  NOR3_X4 U3256 ( .A1(n2029), .A2(n2030), .A3(n2166), .ZN(n2039) );
  NAND2_X2 U3257 ( .A1(n2319), .A2(n2032), .ZN(n2033) );
  INV_X4 U3258 ( .A(n2166), .ZN(n2031) );
  NOR2_X4 U3259 ( .A1(n2031), .A2(n2033), .ZN(n2037) );
  NOR2_X4 U3260 ( .A1(n2038), .A2(n2039), .ZN(n2110) );
  INV_X4 U3261 ( .A(n2040), .ZN(n2042) );
  XNOR2_X2 U3262 ( .A(n2047), .B(n2052), .ZN(n2048) );
  OAI21_X4 U3263 ( .B1(n973), .B2(n2051), .A(net154699), .ZN(n2136) );
  INV_X4 U3264 ( .A(x[21]), .ZN(n2052) );
  INV_X4 U3265 ( .A(x[22]), .ZN(n2057) );
  NOR2_X4 U3266 ( .A1(x[22]), .A2(x[21]), .ZN(n2054) );
  INV_X4 U3267 ( .A(n2122), .ZN(n2055) );
  NAND2_X2 U3268 ( .A1(x[20]), .A2(net153769), .ZN(n2058) );
  INV_X4 U3269 ( .A(net154623), .ZN(net154721) );
  XNOR2_X2 U3270 ( .A(n2136), .B(n2135), .ZN(net154667) );
  NAND2_X2 U3271 ( .A1(x[19]), .A2(n1183), .ZN(n2059) );
  XNOR2_X2 U3272 ( .A(net156803), .B(n2159), .ZN(n2060) );
  XNOR2_X2 U3273 ( .A(n2061), .B(n2060), .ZN(net154349) );
  INV_X4 U3274 ( .A(n2080), .ZN(n2063) );
  NAND2_X2 U3275 ( .A1(n2134), .A2(n2064), .ZN(n2069) );
  INV_X4 U3276 ( .A(n2065), .ZN(n2081) );
  AOI221_X2 U3277 ( .B1(n2081), .B2(n2080), .C1(net154288), .C2(n2067), .A(
        net154711), .ZN(n2068) );
  NAND2_X2 U3278 ( .A1(n2103), .A2(n2170), .ZN(n2073) );
  NAND2_X2 U3279 ( .A1(n2103), .A2(net153937), .ZN(n2072) );
  XNOR2_X2 U3280 ( .A(n2076), .B(net157532), .ZN(net154622) );
  NAND2_X2 U3281 ( .A1(n2084), .A2(n2083), .ZN(n2239) );
  INV_X4 U3282 ( .A(x[23]), .ZN(n2089) );
  INV_X4 U3283 ( .A(x[23]), .ZN(n2121) );
  XNOR2_X2 U3284 ( .A(n2596), .B(n2121), .ZN(n2088) );
  NAND2_X2 U3285 ( .A1(x[21]), .A2(net153769), .ZN(n2090) );
  INV_X4 U3286 ( .A(n2140), .ZN(n2091) );
  NAND2_X2 U3287 ( .A1(x[20]), .A2(n1183), .ZN(n2092) );
  INV_X4 U3288 ( .A(n2273), .ZN(n2094) );
  XNOR2_X2 U3289 ( .A(net156296), .B(n2094), .ZN(n2322) );
  INV_X4 U3290 ( .A(n2097), .ZN(n2100) );
  INV_X4 U3291 ( .A(n2325), .ZN(n2174) );
  NAND2_X2 U3292 ( .A1(n2104), .A2(n2105), .ZN(n2106) );
  NAND2_X2 U3293 ( .A1(n2106), .A2(n2170), .ZN(n2109) );
  NAND2_X2 U3294 ( .A1(n2107), .A2(n2106), .ZN(n2108) );
  NAND2_X2 U3295 ( .A1(x[21]), .A2(n1183), .ZN(n2111) );
  NOR2_X4 U3296 ( .A1(n642), .A2(n2117), .ZN(n2119) );
  INV_X4 U3297 ( .A(x[24]), .ZN(n2120) );
  NAND3_X4 U3298 ( .A1(net154629), .A2(n1181), .A3(n2123), .ZN(n2228) );
  NAND2_X2 U3299 ( .A1(x[24]), .A2(n2606), .ZN(n2124) );
  NAND2_X2 U3300 ( .A1(x[22]), .A2(net153769), .ZN(n2126) );
  XNOR2_X2 U3301 ( .A(n2133), .B(n1003), .ZN(n2141) );
  NAND2_X2 U3302 ( .A1(net154038), .A2(n2521), .ZN(n2149) );
  XNOR2_X2 U3303 ( .A(n2136), .B(n2135), .ZN(net154291) );
  INV_X4 U3304 ( .A(n2137), .ZN(n2148) );
  NOR3_X4 U3305 ( .A1(net154595), .A2(n2147), .A3(net154588), .ZN(n2143) );
  NAND3_X2 U3306 ( .A1(n533), .A2(n2142), .A3(net154341), .ZN(n2162) );
  INV_X4 U3307 ( .A(n2159), .ZN(n2157) );
  INV_X4 U3308 ( .A(n2322), .ZN(n2303) );
  NAND2_X2 U3309 ( .A1(n2308), .A2(n2177), .ZN(n2175) );
  NAND4_X2 U3310 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2170), .ZN(n2184)
         );
  NOR4_X2 U3311 ( .A1(n2180), .A2(n2567), .A3(n2179), .A4(n2178), .ZN(n2181)
         );
  NOR3_X4 U3312 ( .A1(n2186), .A2(net156296), .A3(net154031), .ZN(n2330) );
  NAND2_X2 U3313 ( .A1(x[25]), .A2(n2606), .ZN(n2235) );
  INV_X4 U3314 ( .A(x[25]), .ZN(n2191) );
  XNOR2_X2 U3315 ( .A(n2228), .B(n2191), .ZN(n2231) );
  NAND2_X2 U3316 ( .A1(x[24]), .A2(net155884), .ZN(n2192) );
  XNOR2_X2 U3317 ( .A(n2195), .B(n2194), .ZN(n2232) );
  INV_X4 U3318 ( .A(n2196), .ZN(n2334) );
  INV_X4 U3319 ( .A(n2202), .ZN(n2242) );
  INV_X4 U3320 ( .A(n2239), .ZN(n2200) );
  NOR2_X4 U3321 ( .A1(n2242), .A2(n2200), .ZN(n2201) );
  NAND3_X4 U3322 ( .A1(n2207), .A2(net157532), .A3(net154499), .ZN(n2363) );
  XNOR2_X2 U3323 ( .A(n2333), .B(n2334), .ZN(n2506) );
  NAND2_X2 U3324 ( .A1(x[22]), .A2(n1183), .ZN(n2211) );
  INV_X4 U3325 ( .A(n2552), .ZN(n2546) );
  XNOR2_X2 U3326 ( .A(n880), .B(n2546), .ZN(n2263) );
  XNOR2_X2 U3327 ( .A(n2264), .B(n2263), .ZN(net153696) );
  XNOR2_X2 U3328 ( .A(n2213), .B(n553), .ZN(result[25]) );
  INV_X4 U3329 ( .A(n2214), .ZN(n2215) );
  NAND3_X4 U3330 ( .A1(n2220), .A2(n2221), .A3(n538), .ZN(n2223) );
  NAND2_X2 U3331 ( .A1(x[24]), .A2(net153769), .ZN(n2227) );
  OAI21_X4 U3332 ( .B1(net155839), .B2(n2375), .A(n2227), .ZN(net154055) );
  INV_X4 U3333 ( .A(n2231), .ZN(n2414) );
  OAI22_X2 U3334 ( .A1(net155885), .A2(n2191), .B1(n2414), .B2(net155857), 
        .ZN(n2367) );
  NAND4_X2 U3335 ( .A1(n1094), .A2(net154616), .A3(n2233), .A4(net154459), 
        .ZN(net154323) );
  OAI21_X4 U3336 ( .B1(n2414), .B2(net155869), .A(n2235), .ZN(n2237) );
  INV_X4 U3337 ( .A(n2407), .ZN(n2370) );
  OAI21_X4 U3338 ( .B1(n2238), .B2(n1176), .A(n2370), .ZN(n2248) );
  NAND2_X2 U3339 ( .A1(n2371), .A2(n2239), .ZN(n2243) );
  INV_X4 U3340 ( .A(n2240), .ZN(n2241) );
  NAND2_X2 U3341 ( .A1(x[23]), .A2(n1183), .ZN(n2249) );
  INV_X4 U3342 ( .A(net153986), .ZN(net154438) );
  XNOR2_X2 U3343 ( .A(net153829), .B(net154438), .ZN(n2563) );
  INV_X4 U3344 ( .A(net154143), .ZN(net153550) );
  INV_X4 U3345 ( .A(n2269), .ZN(n2251) );
  XNOR2_X2 U3346 ( .A(n2254), .B(n619), .ZN(n2262) );
  XOR2_X2 U3347 ( .A(n2256), .B(n2255), .Z(n2261) );
  XNOR2_X2 U3348 ( .A(n2264), .B(n2263), .ZN(n2565) );
  AOI21_X4 U3349 ( .B1(n2275), .B2(n584), .A(n2306), .ZN(n2297) );
  NAND2_X2 U3350 ( .A1(n2279), .A2(n2277), .ZN(n2281) );
  NAND2_X2 U3351 ( .A1(n2283), .A2(n2282), .ZN(n2285) );
  NAND3_X4 U3352 ( .A1(n2297), .A2(n2296), .A3(n2295), .ZN(net153700) );
  XNOR2_X2 U3353 ( .A(n2303), .B(n2323), .ZN(n2304) );
  OAI21_X4 U3354 ( .B1(n2304), .B2(n2305), .A(net153533), .ZN(net153936) );
  INV_X4 U3355 ( .A(n2307), .ZN(n2327) );
  OAI21_X4 U3356 ( .B1(net155985), .B2(n2311), .A(n883), .ZN(n2312) );
  OAI21_X4 U3357 ( .B1(n2313), .B2(n2314), .A(n2312), .ZN(n2315) );
  XNOR2_X2 U3358 ( .A(n2317), .B(net153550), .ZN(result[26]) );
  INV_X4 U3359 ( .A(n2318), .ZN(n2426) );
  NAND2_X2 U3360 ( .A1(net154423), .A2(n596), .ZN(n2321) );
  NAND2_X2 U3361 ( .A1(n2872), .A2(net153533), .ZN(n2436) );
  OAI21_X2 U3362 ( .B1(n2436), .B2(n2328), .A(n586), .ZN(n2331) );
  NAND2_X2 U3363 ( .A1(net154322), .A2(net154323), .ZN(n2332) );
  XNOR2_X2 U3364 ( .A(n2332), .B(net158084), .ZN(n2508) );
  XNOR2_X2 U3365 ( .A(n2333), .B(n2334), .ZN(n2665) );
  INV_X4 U3366 ( .A(n2335), .ZN(n2338) );
  NOR2_X4 U3367 ( .A1(n2347), .A2(n2342), .ZN(n2343) );
  NAND2_X2 U3368 ( .A1(net158099), .A2(net154091), .ZN(n2351) );
  NAND2_X2 U3369 ( .A1(net154280), .A2(n2354), .ZN(n2355) );
  AOI211_X4 U3370 ( .C1(n2355), .C2(n2356), .A(n1095), .B(n840), .ZN(net154277) );
  NAND4_X2 U3371 ( .A1(net157527), .A2(net157773), .A3(net158305), .A4(
        net158099), .ZN(n2573) );
  INV_X4 U3372 ( .A(x[27]), .ZN(n2361) );
  NAND2_X2 U3373 ( .A1(x[27]), .A2(n2358), .ZN(n2360) );
  INV_X4 U3374 ( .A(x[26]), .ZN(n2362) );
  OAI22_X2 U3375 ( .A1(net155896), .A2(n2191), .B1(n2414), .B2(net155841), 
        .ZN(net154234) );
  INV_X4 U3376 ( .A(n2409), .ZN(n2368) );
  NAND2_X2 U3377 ( .A1(n2381), .A2(n2409), .ZN(n2373) );
  INV_X4 U3378 ( .A(x[24]), .ZN(n2376) );
  OAI22_X2 U3379 ( .A1(n2705), .A2(n2376), .B1(net155827), .B2(n2375), .ZN(
        net153953) );
  INV_X4 U3380 ( .A(net153953), .ZN(net154244) );
  XNOR2_X2 U3381 ( .A(net154083), .B(net154244), .ZN(n2576) );
  INV_X4 U3382 ( .A(n2454), .ZN(n2380) );
  XNOR2_X2 U3383 ( .A(n2383), .B(net154117), .ZN(n2384) );
  INV_X4 U3384 ( .A(n2430), .ZN(n2395) );
  INV_X4 U3385 ( .A(n2505), .ZN(n2392) );
  NOR2_X4 U3386 ( .A1(n2392), .A2(net153876), .ZN(n2393) );
  NAND3_X2 U3387 ( .A1(n2449), .A2(net154127), .A3(n2428), .ZN(n2397) );
  NAND2_X2 U3388 ( .A1(x[28]), .A2(n2399), .ZN(n2401) );
  OAI22_X2 U3389 ( .A1(net155885), .A2(n2361), .B1(net155855), .B2(n2542), 
        .ZN(n2460) );
  INV_X4 U3390 ( .A(n2460), .ZN(n2402) );
  XNOR2_X2 U3391 ( .A(n2403), .B(n2402), .ZN(n2610) );
  INV_X4 U3392 ( .A(n2610), .ZN(n2458) );
  XNOR2_X2 U3393 ( .A(n2458), .B(n2444), .ZN(n2412) );
  OAI21_X4 U3394 ( .B1(net154205), .B2(n916), .A(n2409), .ZN(n2404) );
  NAND2_X2 U3395 ( .A1(x[25]), .A2(n1183), .ZN(n2413) );
  INV_X4 U3396 ( .A(n2571), .ZN(n2415) );
  XNOR2_X2 U3397 ( .A(n606), .B(n2415), .ZN(n2578) );
  INV_X4 U3398 ( .A(n2416), .ZN(n2493) );
  OAI21_X2 U3399 ( .B1(n2436), .B2(n2421), .A(n2420), .ZN(n2423) );
  XNOR2_X2 U3400 ( .A(n2424), .B(n2493), .ZN(result[28]) );
  INV_X4 U3401 ( .A(n2427), .ZN(n2494) );
  INV_X4 U3402 ( .A(net154151), .ZN(net153621) );
  NAND3_X2 U3403 ( .A1(net158305), .A2(n2516), .A3(net157527), .ZN(n2482) );
  OAI211_X2 U3404 ( .C1(n2436), .C2(n2328), .A(n586), .B(n2438), .ZN(n2441) );
  INV_X4 U3405 ( .A(n2450), .ZN(n2447) );
  NAND3_X2 U3406 ( .A1(n2449), .A2(net154127), .A3(n2448), .ZN(n2453) );
  AOI21_X2 U3407 ( .B1(n2486), .B2(net158270), .A(net154083), .ZN(n2451) );
  NAND2_X2 U3408 ( .A1(n2717), .A2(n2499), .ZN(n2483) );
  OAI21_X4 U3409 ( .B1(n2540), .B2(n2539), .A(n2615), .ZN(n2501) );
  INV_X4 U3410 ( .A(x[28]), .ZN(n2461) );
  INV_X4 U3411 ( .A(x[29]), .ZN(n2469) );
  INV_X4 U3412 ( .A(x[29]), .ZN(n2467) );
  NOR2_X4 U3413 ( .A1(x[26]), .A2(n2600), .ZN(n2466) );
  NOR2_X4 U3414 ( .A1(x[28]), .A2(x[27]), .ZN(n2463) );
  NAND2_X2 U3415 ( .A1(n2463), .A2(n2467), .ZN(n2597) );
  NOR2_X4 U3416 ( .A1(x[25]), .A2(n2597), .ZN(n2464) );
  NAND3_X4 U3417 ( .A1(n2466), .A2(n2465), .A3(n2464), .ZN(n2529) );
  OAI21_X4 U3418 ( .B1(n2468), .B2(n2467), .A(n2529), .ZN(n2686) );
  OAI22_X2 U3419 ( .A1(net155896), .A2(n2361), .B1(net155839), .B2(n2542), 
        .ZN(n2502) );
  XNOR2_X2 U3420 ( .A(n2616), .B(n2502), .ZN(n2470) );
  XNOR2_X2 U3421 ( .A(n2501), .B(n2470), .ZN(n2627) );
  NAND2_X2 U3422 ( .A1(x[26]), .A2(n1183), .ZN(n2471) );
  INV_X4 U3423 ( .A(n2581), .ZN(n2473) );
  XNOR2_X2 U3424 ( .A(n2649), .B(n2473), .ZN(n2474) );
  NAND2_X2 U3425 ( .A1(net156089), .A2(n2484), .ZN(n2480) );
  NAND3_X2 U3426 ( .A1(n1082), .A2(net154295), .A3(n2481), .ZN(n2491) );
  AOI21_X4 U3427 ( .B1(n2487), .B2(net154083), .A(n2485), .ZN(n2489) );
  NAND3_X2 U3428 ( .A1(n2487), .A2(n2486), .A3(net158270), .ZN(n2488) );
  AOI22_X2 U3429 ( .A1(n2496), .A2(net158256), .B1(net153550), .B2(n2495), 
        .ZN(n2497) );
  AOI21_X4 U3430 ( .B1(n2649), .B2(n2504), .A(n2650), .ZN(n2805) );
  NAND3_X2 U3431 ( .A1(n1169), .A2(net153829), .A3(net153831), .ZN(n2633) );
  NAND3_X4 U3432 ( .A1(n2478), .A2(n2813), .A3(n2516), .ZN(n2723) );
  INV_X4 U3433 ( .A(n2519), .ZN(n2817) );
  OAI211_X2 U3434 ( .C1(n730), .C2(n2521), .A(n2520), .B(net154038), .ZN(
        net154034) );
  NAND2_X2 U3435 ( .A1(x[28]), .A2(net153769), .ZN(n2528) );
  OAI21_X4 U3436 ( .B1(net155839), .B2(n2594), .A(n2528), .ZN(n2625) );
  INV_X4 U3437 ( .A(x[30]), .ZN(n2532) );
  XNOR2_X2 U3438 ( .A(x[30]), .B(n2530), .ZN(n2531) );
  INV_X4 U3439 ( .A(n2531), .ZN(n2704) );
  XNOR2_X2 U3440 ( .A(n2618), .B(n565), .ZN(n2678) );
  XNOR2_X2 U3441 ( .A(n2678), .B(n2625), .ZN(net154006) );
  INV_X4 U3442 ( .A(n2614), .ZN(n2537) );
  INV_X4 U3443 ( .A(n2615), .ZN(n2536) );
  OAI21_X4 U3444 ( .B1(n2540), .B2(n2539), .A(n2538), .ZN(n2621) );
  NAND2_X2 U3445 ( .A1(x[27]), .A2(n1183), .ZN(n2541) );
  INV_X4 U3446 ( .A(net154001), .ZN(net153930) );
  NOR2_X4 U3447 ( .A1(n2545), .A2(n2546), .ZN(n2557) );
  AOI21_X4 U3448 ( .B1(n1084), .B2(n1002), .A(n2558), .ZN(n2554) );
  NAND2_X2 U3449 ( .A1(n2552), .A2(n2518), .ZN(n2560) );
  AOI21_X4 U3450 ( .B1(n1084), .B2(n2559), .A(n2558), .ZN(n2561) );
  XNOR2_X2 U3451 ( .A(n2562), .B(net153975), .ZN(n2589) );
  XNOR2_X2 U3452 ( .A(n2564), .B(n2563), .ZN(net153545) );
  NOR2_X4 U3453 ( .A1(n2566), .A2(n2567), .ZN(net153960) );
  AOI21_X4 U3454 ( .B1(net153958), .B2(net153700), .A(net153959), .ZN(n2570)
         );
  INV_X4 U3455 ( .A(n2573), .ZN(n2574) );
  XNOR2_X2 U3456 ( .A(n2577), .B(n2576), .ZN(n2580) );
  XNOR2_X2 U3457 ( .A(n2579), .B(n2578), .ZN(n2863) );
  OAI21_X4 U3458 ( .B1(net153942), .B2(n2580), .A(n2863), .ZN(n2583) );
  NAND3_X4 U3459 ( .A1(n2583), .A2(n686), .A3(n2729), .ZN(n2689) );
  INV_X4 U3460 ( .A(net153788), .ZN(net153598) );
  NAND2_X2 U3461 ( .A1(n2591), .A2(n2590), .ZN(n2593) );
  OAI22_X2 U3462 ( .A1(n2705), .A2(n2461), .B1(net155827), .B2(n2594), .ZN(
        n2695) );
  INV_X4 U3463 ( .A(n2695), .ZN(n2748) );
  NAND2_X2 U3464 ( .A1(x[29]), .A2(net153769), .ZN(n2595) );
  INV_X4 U3465 ( .A(n2657), .ZN(n2620) );
  INV_X4 U3466 ( .A(n2597), .ZN(n2602) );
  INV_X4 U3467 ( .A(n2598), .ZN(n2599) );
  NAND4_X2 U3468 ( .A1(n2465), .A2(n2532), .A3(n2602), .A4(n2601), .ZN(n2604)
         );
  INV_X4 U3469 ( .A(x[31]), .ZN(n2603) );
  XNOR2_X2 U3470 ( .A(n2604), .B(n2603), .ZN(n2605) );
  INV_X4 U3471 ( .A(n2605), .ZN(n2804) );
  NAND2_X2 U3472 ( .A1(x[31]), .A2(n2606), .ZN(n2607) );
  OAI21_X4 U3473 ( .B1(n2804), .B2(net155869), .A(n2607), .ZN(n2707) );
  INV_X4 U3474 ( .A(n2707), .ZN(n2674) );
  OAI22_X2 U3475 ( .A1(net155885), .A2(n2532), .B1(n2704), .B2(net155857), 
        .ZN(n2675) );
  INV_X4 U3476 ( .A(n2675), .ZN(n2608) );
  XNOR2_X2 U3477 ( .A(n2674), .B(n2608), .ZN(n2800) );
  INV_X4 U3478 ( .A(n2800), .ZN(n2786) );
  NOR2_X4 U3479 ( .A1(n2613), .A2(n2677), .ZN(n2617) );
  OAI21_X4 U3480 ( .B1(n2616), .B2(n2615), .A(n2614), .ZN(n2676) );
  NAND2_X2 U3481 ( .A1(n2618), .A2(n565), .ZN(n2783) );
  XNOR2_X2 U3482 ( .A(n2786), .B(n2653), .ZN(n2652) );
  XNOR2_X2 U3483 ( .A(n1080), .B(n2748), .ZN(n2826) );
  XNOR2_X2 U3484 ( .A(n2623), .B(n850), .ZN(n2624) );
  INV_X4 U3485 ( .A(net153863), .ZN(net153881) );
  NAND3_X4 U3486 ( .A1(n1167), .A2(n818), .A3(net158266), .ZN(n2642) );
  OAI21_X4 U3487 ( .B1(n2637), .B2(n2636), .A(n2635), .ZN(n2638) );
  XNOR2_X2 U3488 ( .A(n2826), .B(n2694), .ZN(n2749) );
  XNOR2_X2 U3489 ( .A(n2786), .B(n2657), .ZN(n2647) );
  NOR2_X4 U3490 ( .A1(n2650), .A2(n2649), .ZN(n2651) );
  XNOR2_X2 U3491 ( .A(n2786), .B(n2653), .ZN(n2656) );
  INV_X4 U3492 ( .A(n2658), .ZN(n2659) );
  INV_X4 U3493 ( .A(n2667), .ZN(n2668) );
  OAI21_X4 U3494 ( .B1(net153823), .B2(n2669), .A(n2668), .ZN(n2811) );
  NAND2_X2 U3495 ( .A1(n2741), .A2(n2743), .ZN(n2688) );
  NAND2_X2 U3496 ( .A1(x[30]), .A2(net153769), .ZN(n2672) );
  OAI22_X2 U3497 ( .A1(n2603), .A2(net155885), .B1(n2804), .B2(net155855), 
        .ZN(n2708) );
  INV_X4 U3498 ( .A(n2708), .ZN(n2673) );
  XNOR2_X2 U3499 ( .A(n2674), .B(n2673), .ZN(n2714) );
  XNOR2_X2 U3500 ( .A(n2715), .B(n2714), .ZN(n2684) );
  NAND2_X2 U3501 ( .A1(n2675), .A2(n2707), .ZN(n2798) );
  NAND2_X2 U3502 ( .A1(n2800), .A2(n2798), .ZN(n2681) );
  XNOR2_X2 U3503 ( .A(n2684), .B(n2716), .ZN(n2789) );
  NAND2_X2 U3504 ( .A1(x[29]), .A2(n1183), .ZN(n2685) );
  INV_X4 U3505 ( .A(n2830), .ZN(n2687) );
  XNOR2_X2 U3506 ( .A(n2895), .B(n2687), .ZN(n2744) );
  XNOR2_X2 U3507 ( .A(n2688), .B(n2744), .ZN(n2731) );
  INV_X4 U3508 ( .A(n2731), .ZN(n2750) );
  INV_X4 U3509 ( .A(n1022), .ZN(n2690) );
  OAI22_X2 U3510 ( .A1(n2705), .A2(n2532), .B1(n2704), .B2(net155835), .ZN(
        n2776) );
  NAND2_X2 U3511 ( .A1(net153769), .A2(x[31]), .ZN(n2706) );
  NAND2_X2 U3512 ( .A1(n2708), .A2(n2707), .ZN(n2910) );
  NAND2_X2 U3513 ( .A1(n2714), .A2(n2910), .ZN(n2802) );
  NAND2_X2 U3514 ( .A1(n2802), .A2(n2798), .ZN(n2781) );
  INV_X4 U3515 ( .A(n2910), .ZN(n2710) );
  INV_X4 U3516 ( .A(n2714), .ZN(n2909) );
  NAND2_X2 U3517 ( .A1(n2890), .A2(n2894), .ZN(n2773) );
  NAND2_X2 U3518 ( .A1(n2895), .A2(n2894), .ZN(n2772) );
  INV_X4 U3519 ( .A(n2719), .ZN(n2807) );
  NAND3_X2 U3520 ( .A1(n1123), .A2(n2723), .A3(n2722), .ZN(n2739) );
  XNOR2_X2 U3521 ( .A(n2726), .B(n2727), .ZN(n2877) );
  INV_X4 U3522 ( .A(n2728), .ZN(n2730) );
  NAND2_X2 U3523 ( .A1(n756), .A2(n2736), .ZN(n2737) );
  XNOR2_X2 U3524 ( .A(n2742), .B(n1060), .ZN(n2763) );
  NAND2_X2 U3525 ( .A1(n2741), .A2(n2743), .ZN(n2745) );
  NOR3_X4 U3526 ( .A1(n2747), .A2(n2834), .A3(n2748), .ZN(n2780) );
  INV_X4 U3527 ( .A(n2752), .ZN(n2754) );
  OAI21_X4 U3528 ( .B1(n2759), .B2(n2758), .A(n2757), .ZN(n2760) );
  INV_X4 U3529 ( .A(n2764), .ZN(n2765) );
  OAI21_X4 U3530 ( .B1(n2779), .B2(n705), .A(n2778), .ZN(net153667) );
  INV_X4 U3531 ( .A(n2908), .ZN(n2782) );
  NOR2_X4 U3532 ( .A1(n2782), .A2(n2781), .ZN(n2788) );
  NAND3_X2 U3533 ( .A1(n2785), .A2(n2784), .A3(n2783), .ZN(n2797) );
  NAND2_X2 U3534 ( .A1(n2894), .A2(n2898), .ZN(n2790) );
  NAND2_X2 U3535 ( .A1(n2794), .A2(n2793), .ZN(n2795) );
  OAI21_X4 U3536 ( .B1(n2796), .B2(n2829), .A(n2795), .ZN(net153525) );
  INV_X4 U3537 ( .A(n2801), .ZN(n2911) );
  XNOR2_X2 U3538 ( .A(n2902), .B(n2908), .ZN(n2845) );
  NAND2_X2 U3539 ( .A1(n1183), .A2(x[31]), .ZN(n2803) );
  XNOR2_X2 U3540 ( .A(n2845), .B(n2907), .ZN(net153526) );
  INV_X4 U3541 ( .A(net153517), .ZN(net153600) );
  INV_X4 U3542 ( .A(n2812), .ZN(n2824) );
  NOR2_X4 U3543 ( .A1(n656), .A2(n2816), .ZN(n2820) );
  OAI21_X4 U3544 ( .B1(n2823), .B2(n2822), .A(n2821), .ZN(n2847) );
  XNOR2_X2 U3545 ( .A(n2826), .B(n2825), .ZN(n2879) );
  NAND2_X2 U3546 ( .A1(net153600), .A2(n2879), .ZN(n2827) );
  INV_X4 U3547 ( .A(n2827), .ZN(n2837) );
  NOR2_X4 U3548 ( .A1(n2837), .A2(net153598), .ZN(n2840) );
  NAND2_X2 U3549 ( .A1(n2830), .A2(n2895), .ZN(n2831) );
  XNOR2_X2 U3550 ( .A(n2832), .B(n2831), .ZN(n2833) );
  NOR2_X4 U3551 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  NOR3_X4 U3552 ( .A1(n2839), .A2(n2840), .A3(n2882), .ZN(n2862) );
  NAND3_X2 U3553 ( .A1(n1052), .A2(n2851), .A3(n2850), .ZN(n2852) );
  OAI21_X4 U3554 ( .B1(n2853), .B2(n2854), .A(n2852), .ZN(n2855) );
  AOI21_X4 U3555 ( .B1(net153559), .B2(net156776), .A(net153561), .ZN(n2860)
         );
  NAND3_X2 U3556 ( .A1(n2870), .A2(net153548), .A3(net153549), .ZN(n2871) );
  NAND3_X2 U3557 ( .A1(n2868), .A2(n2869), .A3(n2870), .ZN(n2873) );
  NAND2_X2 U3558 ( .A1(n2874), .A2(n2873), .ZN(n2886) );
  NOR2_X4 U3559 ( .A1(n2838), .A2(n2881), .ZN(n2883) );
  INV_X4 U3560 ( .A(n2898), .ZN(n2899) );
  NAND2_X2 U3561 ( .A1(n2903), .A2(n2908), .ZN(n2904) );
  OAI21_X4 U3562 ( .B1(n2906), .B2(n2905), .A(n2904), .ZN(n2916) );
  INV_X4 U3563 ( .A(n2907), .ZN(n2914) );
  XNOR2_X2 U3564 ( .A(n2909), .B(n2908), .ZN(n2913) );
  NAND2_X2 U3565 ( .A1(n2911), .A2(n2910), .ZN(n2912) );
  FA_X1 U3566 ( .A(n2914), .B(n2913), .CI(n2912), .S(n2915) );
  XNOR2_X2 U3567 ( .A(n2916), .B(n2915), .ZN(n2917) );
endmodule

