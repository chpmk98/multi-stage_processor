
module pp ( clk, regRst, pcIn, pcRst, iaddr, inst, daddr, drData, dwData, dWr, 
        dSize, dpcHold, difHold, didHold, difKill, didKill, daluKill, didMult, 
        idRegWr, aluRegWrOut, wbBusWh, wbRegWrh, wbRwh, ifInst );
  input [31:0] pcIn;
  output [31:0] iaddr;
  input [31:0] inst;
  output [31:0] daddr;
  input [31:0] drData;
  output [31:0] dwData;
  output [1:0] dSize;
  output [31:0] wbBusWh;
  output [4:0] wbRwh;
  output [31:0] ifInst;
  input clk, regRst, pcRst;
  output dWr, dpcHold, difHold, didHold, difKill, didKill, daluKill, didMult,
         idRegWr, aluRegWrOut, wbRegWrh;
  wire   aluifJRflag, ifOut_95_, ifOut_94_, ifOut_93_, ifOut_92_, ifOut_91_,
         ifOut_90_, ifOut_89_, ifOut_88_, ifOut_87_, ifOut_86_, ifOut_85_,
         ifOut_84_, ifOut_83_, ifOut_82_, ifOut_81_, ifOut_80_, ifOut_79_,
         ifOut_78_, ifOut_77_, ifOut_76_, ifOut_75_, ifOut_74_, ifOut_73_,
         ifOut_72_, ifOut_71_, ifOut_70_, ifOut_69_, ifOut_68_, ifOut_67_,
         ifOut_66_, ifOut_65_, ifOut_64_, ifOut_31_, ifOut_30_, ifOut_29_,
         ifOut_28_, ifOut_27_, ifOut_26_, ifOut_25_, ifOut_24_, ifOut_23_,
         ifOut_22_, ifOut_21_, ifOut_20_, ifOut_19_, ifOut_18_, ifOut_17_,
         ifOut_16_, ifOut_15_, ifOut_14_, ifOut_13_, ifOut_12_, ifOut_11_,
         ifOut_10_, ifOut_9_, ifOut_8_, ifOut_7_, ifOut_6_, ifOut_5_, ifOut_4_,
         ifOut_3_, ifOut_2_, ifOut_1_, ifOut_0_, idOut_117_, idOut_116_,
         idOut_115_, idOut_114_, idOut_113_, idOut_112_, idOut_111_,
         idOut_110_, idOut_109_, idOut_108_, idOut_107_, idOut_106_,
         idOut_105_, idOut_104_, idOut_103_, idOut_102_, idOut_101_,
         idOut_100_, idOut_99_, idOut_98_, idOut_97_, idOut_96_, idOut_95_,
         idOut_94_, idOut_93_, idOut_92_, idOut_91_, idOut_90_, idOut_89_,
         idOut_88_, idOut_87_, idOut_86_, idOut_75_, idOut_74_, idOut_73_,
         idOut_72_, idOut_71_, idOut_70_, idOut_69_, idOut_68_, idOut_67_,
         idOut_66_, idOut_65_, idOut_64_, idOut_63_, idOut_62_, idOut_61_,
         idOut_60_, idOut_59_, idOut_58_, idOut_57_, idOut_56_, idOut_55_,
         idOut_54_, idOut_53_, idOut_52_, idOut_51_, idOut_50_, idOut_49_,
         idOut_48_, idOut_47_, idOut_46_, idOut_45_, idOut_44_, idOut_43_,
         idOut_42_, idOut_41_, idOut_40_, idOut_39_, idOut_38_, idOut_34_,
         idOut_33_, idOut_32_, idOut_31_, idOut_29_, idOut_28_, idOut_26_,
         idOut_25_, idOut_24_, idOut_23_, idOut_22_, idOut_21_, idOut_20_,
         idOut_19_, idOut_18_, idOut_17_, idOut_16_, difHold, aluDExtOp,
         aluJAL, aluMem2Reg, MoLanBoJ, idBoi_temPC_0_, idBoi_temPC_1_,
         idBoi_temPC_2_, regBoiz_regfile_31__31_, regBoiz_regfile_31__30_,
         regBoiz_regfile_31__29_, regBoiz_regfile_31__28_,
         regBoiz_regfile_31__27_, regBoiz_regfile_31__26_,
         regBoiz_regfile_31__25_, regBoiz_regfile_31__24_,
         regBoiz_regfile_31__23_, regBoiz_regfile_31__22_,
         regBoiz_regfile_31__21_, regBoiz_regfile_31__20_,
         regBoiz_regfile_31__19_, regBoiz_regfile_31__18_,
         regBoiz_regfile_31__17_, regBoiz_regfile_31__16_,
         regBoiz_regfile_31__15_, regBoiz_regfile_31__14_,
         regBoiz_regfile_31__13_, regBoiz_regfile_31__12_,
         regBoiz_regfile_31__11_, regBoiz_regfile_31__10_,
         regBoiz_regfile_31__9_, regBoiz_regfile_31__8_,
         regBoiz_regfile_31__7_, regBoiz_regfile_31__6_,
         regBoiz_regfile_31__5_, regBoiz_regfile_31__4_,
         regBoiz_regfile_31__3_, regBoiz_regfile_31__2_,
         regBoiz_regfile_31__1_, regBoiz_regfile_31__0_,
         regBoiz_regfile_30__31_, regBoiz_regfile_30__30_,
         regBoiz_regfile_30__29_, regBoiz_regfile_30__28_,
         regBoiz_regfile_30__27_, regBoiz_regfile_30__26_,
         regBoiz_regfile_30__25_, regBoiz_regfile_30__24_,
         regBoiz_regfile_30__23_, regBoiz_regfile_30__22_,
         regBoiz_regfile_30__21_, regBoiz_regfile_30__20_,
         regBoiz_regfile_30__19_, regBoiz_regfile_30__18_,
         regBoiz_regfile_30__17_, regBoiz_regfile_30__16_,
         regBoiz_regfile_30__15_, regBoiz_regfile_30__14_,
         regBoiz_regfile_30__13_, regBoiz_regfile_30__12_,
         regBoiz_regfile_30__11_, regBoiz_regfile_30__10_,
         regBoiz_regfile_30__9_, regBoiz_regfile_30__8_,
         regBoiz_regfile_30__7_, regBoiz_regfile_30__6_,
         regBoiz_regfile_30__5_, regBoiz_regfile_30__4_,
         regBoiz_regfile_30__3_, regBoiz_regfile_30__2_,
         regBoiz_regfile_30__1_, regBoiz_regfile_30__0_,
         regBoiz_regfile_29__31_, regBoiz_regfile_29__30_,
         regBoiz_regfile_29__29_, regBoiz_regfile_29__28_,
         regBoiz_regfile_29__27_, regBoiz_regfile_29__26_,
         regBoiz_regfile_29__25_, regBoiz_regfile_29__24_,
         regBoiz_regfile_29__23_, regBoiz_regfile_29__22_,
         regBoiz_regfile_29__21_, regBoiz_regfile_29__20_,
         regBoiz_regfile_29__19_, regBoiz_regfile_29__18_,
         regBoiz_regfile_29__17_, regBoiz_regfile_29__16_,
         regBoiz_regfile_29__15_, regBoiz_regfile_29__14_,
         regBoiz_regfile_29__13_, regBoiz_regfile_29__12_,
         regBoiz_regfile_29__11_, regBoiz_regfile_29__10_,
         regBoiz_regfile_29__9_, regBoiz_regfile_29__8_,
         regBoiz_regfile_29__7_, regBoiz_regfile_29__6_,
         regBoiz_regfile_29__5_, regBoiz_regfile_29__4_,
         regBoiz_regfile_29__3_, regBoiz_regfile_29__2_,
         regBoiz_regfile_29__1_, regBoiz_regfile_29__0_,
         regBoiz_regfile_28__31_, regBoiz_regfile_28__30_,
         regBoiz_regfile_28__29_, regBoiz_regfile_28__28_,
         regBoiz_regfile_28__27_, regBoiz_regfile_28__26_,
         regBoiz_regfile_28__25_, regBoiz_regfile_28__24_,
         regBoiz_regfile_28__23_, regBoiz_regfile_28__22_,
         regBoiz_regfile_28__21_, regBoiz_regfile_28__20_,
         regBoiz_regfile_28__19_, regBoiz_regfile_28__18_,
         regBoiz_regfile_28__17_, regBoiz_regfile_28__16_,
         regBoiz_regfile_28__15_, regBoiz_regfile_28__14_,
         regBoiz_regfile_28__13_, regBoiz_regfile_28__12_,
         regBoiz_regfile_28__11_, regBoiz_regfile_28__10_,
         regBoiz_regfile_28__9_, regBoiz_regfile_28__8_,
         regBoiz_regfile_28__7_, regBoiz_regfile_28__6_,
         regBoiz_regfile_28__5_, regBoiz_regfile_28__4_,
         regBoiz_regfile_28__3_, regBoiz_regfile_28__2_,
         regBoiz_regfile_28__1_, regBoiz_regfile_28__0_,
         regBoiz_regfile_27__31_, regBoiz_regfile_27__30_,
         regBoiz_regfile_27__29_, regBoiz_regfile_27__28_,
         regBoiz_regfile_27__27_, regBoiz_regfile_27__26_,
         regBoiz_regfile_27__25_, regBoiz_regfile_27__24_,
         regBoiz_regfile_27__23_, regBoiz_regfile_27__22_,
         regBoiz_regfile_27__21_, regBoiz_regfile_27__20_,
         regBoiz_regfile_27__19_, regBoiz_regfile_27__18_,
         regBoiz_regfile_27__17_, regBoiz_regfile_27__16_,
         regBoiz_regfile_27__15_, regBoiz_regfile_27__14_,
         regBoiz_regfile_27__13_, regBoiz_regfile_27__12_,
         regBoiz_regfile_27__11_, regBoiz_regfile_27__10_,
         regBoiz_regfile_27__9_, regBoiz_regfile_27__8_,
         regBoiz_regfile_27__7_, regBoiz_regfile_27__6_,
         regBoiz_regfile_27__5_, regBoiz_regfile_27__4_,
         regBoiz_regfile_27__3_, regBoiz_regfile_27__2_,
         regBoiz_regfile_27__1_, regBoiz_regfile_27__0_,
         regBoiz_regfile_26__31_, regBoiz_regfile_26__30_,
         regBoiz_regfile_26__29_, regBoiz_regfile_26__28_,
         regBoiz_regfile_26__27_, regBoiz_regfile_26__26_,
         regBoiz_regfile_26__25_, regBoiz_regfile_26__24_,
         regBoiz_regfile_26__23_, regBoiz_regfile_26__22_,
         regBoiz_regfile_26__21_, regBoiz_regfile_26__20_,
         regBoiz_regfile_26__19_, regBoiz_regfile_26__18_,
         regBoiz_regfile_26__17_, regBoiz_regfile_26__16_,
         regBoiz_regfile_26__15_, regBoiz_regfile_26__14_,
         regBoiz_regfile_26__13_, regBoiz_regfile_26__12_,
         regBoiz_regfile_26__11_, regBoiz_regfile_26__10_,
         regBoiz_regfile_26__9_, regBoiz_regfile_26__8_,
         regBoiz_regfile_26__7_, regBoiz_regfile_26__6_,
         regBoiz_regfile_26__5_, regBoiz_regfile_26__4_,
         regBoiz_regfile_26__3_, regBoiz_regfile_26__2_,
         regBoiz_regfile_26__1_, regBoiz_regfile_26__0_,
         regBoiz_regfile_25__31_, regBoiz_regfile_25__30_,
         regBoiz_regfile_25__29_, regBoiz_regfile_25__28_,
         regBoiz_regfile_25__27_, regBoiz_regfile_25__26_,
         regBoiz_regfile_25__25_, regBoiz_regfile_25__24_,
         regBoiz_regfile_25__23_, regBoiz_regfile_25__22_,
         regBoiz_regfile_25__21_, regBoiz_regfile_25__20_,
         regBoiz_regfile_25__19_, regBoiz_regfile_25__18_,
         regBoiz_regfile_25__17_, regBoiz_regfile_25__16_,
         regBoiz_regfile_25__15_, regBoiz_regfile_25__14_,
         regBoiz_regfile_25__13_, regBoiz_regfile_25__12_,
         regBoiz_regfile_25__11_, regBoiz_regfile_25__10_,
         regBoiz_regfile_25__9_, regBoiz_regfile_25__8_,
         regBoiz_regfile_25__7_, regBoiz_regfile_25__6_,
         regBoiz_regfile_25__5_, regBoiz_regfile_25__4_,
         regBoiz_regfile_25__3_, regBoiz_regfile_25__2_,
         regBoiz_regfile_25__1_, regBoiz_regfile_25__0_,
         regBoiz_regfile_24__31_, regBoiz_regfile_24__30_,
         regBoiz_regfile_24__29_, regBoiz_regfile_24__28_,
         regBoiz_regfile_24__27_, regBoiz_regfile_24__26_,
         regBoiz_regfile_24__25_, regBoiz_regfile_24__24_,
         regBoiz_regfile_24__23_, regBoiz_regfile_24__22_,
         regBoiz_regfile_24__21_, regBoiz_regfile_24__20_,
         regBoiz_regfile_24__19_, regBoiz_regfile_24__18_,
         regBoiz_regfile_24__17_, regBoiz_regfile_24__16_,
         regBoiz_regfile_24__15_, regBoiz_regfile_24__14_,
         regBoiz_regfile_24__13_, regBoiz_regfile_24__12_,
         regBoiz_regfile_24__11_, regBoiz_regfile_24__10_,
         regBoiz_regfile_24__9_, regBoiz_regfile_24__8_,
         regBoiz_regfile_24__7_, regBoiz_regfile_24__6_,
         regBoiz_regfile_24__5_, regBoiz_regfile_24__4_,
         regBoiz_regfile_24__3_, regBoiz_regfile_24__2_,
         regBoiz_regfile_24__1_, regBoiz_regfile_24__0_,
         regBoiz_regfile_23__31_, regBoiz_regfile_23__30_,
         regBoiz_regfile_23__29_, regBoiz_regfile_23__28_,
         regBoiz_regfile_23__27_, regBoiz_regfile_23__26_,
         regBoiz_regfile_23__25_, regBoiz_regfile_23__24_,
         regBoiz_regfile_23__23_, regBoiz_regfile_23__22_,
         regBoiz_regfile_23__21_, regBoiz_regfile_23__20_,
         regBoiz_regfile_23__19_, regBoiz_regfile_23__18_,
         regBoiz_regfile_23__17_, regBoiz_regfile_23__16_,
         regBoiz_regfile_23__15_, regBoiz_regfile_23__14_,
         regBoiz_regfile_23__13_, regBoiz_regfile_23__12_,
         regBoiz_regfile_23__11_, regBoiz_regfile_23__10_,
         regBoiz_regfile_23__9_, regBoiz_regfile_23__8_,
         regBoiz_regfile_23__7_, regBoiz_regfile_23__6_,
         regBoiz_regfile_23__5_, regBoiz_regfile_23__4_,
         regBoiz_regfile_23__3_, regBoiz_regfile_23__2_,
         regBoiz_regfile_23__1_, regBoiz_regfile_23__0_,
         regBoiz_regfile_22__31_, regBoiz_regfile_22__30_,
         regBoiz_regfile_22__29_, regBoiz_regfile_22__28_,
         regBoiz_regfile_22__27_, regBoiz_regfile_22__26_,
         regBoiz_regfile_22__25_, regBoiz_regfile_22__24_,
         regBoiz_regfile_22__23_, regBoiz_regfile_22__22_,
         regBoiz_regfile_22__21_, regBoiz_regfile_22__20_,
         regBoiz_regfile_22__19_, regBoiz_regfile_22__18_,
         regBoiz_regfile_22__17_, regBoiz_regfile_22__16_,
         regBoiz_regfile_22__15_, regBoiz_regfile_22__14_,
         regBoiz_regfile_22__13_, regBoiz_regfile_22__12_,
         regBoiz_regfile_22__11_, regBoiz_regfile_22__10_,
         regBoiz_regfile_22__9_, regBoiz_regfile_22__8_,
         regBoiz_regfile_22__7_, regBoiz_regfile_22__6_,
         regBoiz_regfile_22__5_, regBoiz_regfile_22__4_,
         regBoiz_regfile_22__3_, regBoiz_regfile_22__2_,
         regBoiz_regfile_22__1_, regBoiz_regfile_22__0_,
         regBoiz_regfile_21__31_, regBoiz_regfile_21__30_,
         regBoiz_regfile_21__29_, regBoiz_regfile_21__28_,
         regBoiz_regfile_21__27_, regBoiz_regfile_21__26_,
         regBoiz_regfile_21__25_, regBoiz_regfile_21__24_,
         regBoiz_regfile_21__23_, regBoiz_regfile_21__22_,
         regBoiz_regfile_21__21_, regBoiz_regfile_21__20_,
         regBoiz_regfile_21__19_, regBoiz_regfile_21__18_,
         regBoiz_regfile_21__17_, regBoiz_regfile_21__16_,
         regBoiz_regfile_21__15_, regBoiz_regfile_21__14_,
         regBoiz_regfile_21__13_, regBoiz_regfile_21__12_,
         regBoiz_regfile_21__11_, regBoiz_regfile_21__10_,
         regBoiz_regfile_21__9_, regBoiz_regfile_21__8_,
         regBoiz_regfile_21__7_, regBoiz_regfile_21__6_,
         regBoiz_regfile_21__5_, regBoiz_regfile_21__4_,
         regBoiz_regfile_21__3_, regBoiz_regfile_21__2_,
         regBoiz_regfile_21__1_, regBoiz_regfile_21__0_,
         regBoiz_regfile_20__31_, regBoiz_regfile_20__30_,
         regBoiz_regfile_20__29_, regBoiz_regfile_20__28_,
         regBoiz_regfile_20__27_, regBoiz_regfile_20__26_,
         regBoiz_regfile_20__25_, regBoiz_regfile_20__24_,
         regBoiz_regfile_20__23_, regBoiz_regfile_20__22_,
         regBoiz_regfile_20__21_, regBoiz_regfile_20__20_,
         regBoiz_regfile_20__19_, regBoiz_regfile_20__18_,
         regBoiz_regfile_20__17_, regBoiz_regfile_20__16_,
         regBoiz_regfile_20__15_, regBoiz_regfile_20__14_,
         regBoiz_regfile_20__13_, regBoiz_regfile_20__12_,
         regBoiz_regfile_20__11_, regBoiz_regfile_20__10_,
         regBoiz_regfile_20__9_, regBoiz_regfile_20__8_,
         regBoiz_regfile_20__7_, regBoiz_regfile_20__6_,
         regBoiz_regfile_20__5_, regBoiz_regfile_20__4_,
         regBoiz_regfile_20__3_, regBoiz_regfile_20__2_,
         regBoiz_regfile_20__1_, regBoiz_regfile_20__0_,
         regBoiz_regfile_19__31_, regBoiz_regfile_19__30_,
         regBoiz_regfile_19__29_, regBoiz_regfile_19__28_,
         regBoiz_regfile_19__27_, regBoiz_regfile_19__26_,
         regBoiz_regfile_19__25_, regBoiz_regfile_19__24_,
         regBoiz_regfile_19__23_, regBoiz_regfile_19__22_,
         regBoiz_regfile_19__21_, regBoiz_regfile_19__20_,
         regBoiz_regfile_19__19_, regBoiz_regfile_19__18_,
         regBoiz_regfile_19__17_, regBoiz_regfile_19__16_,
         regBoiz_regfile_19__15_, regBoiz_regfile_19__14_,
         regBoiz_regfile_19__13_, regBoiz_regfile_19__12_,
         regBoiz_regfile_19__11_, regBoiz_regfile_19__10_,
         regBoiz_regfile_19__9_, regBoiz_regfile_19__8_,
         regBoiz_regfile_19__7_, regBoiz_regfile_19__6_,
         regBoiz_regfile_19__5_, regBoiz_regfile_19__4_,
         regBoiz_regfile_19__3_, regBoiz_regfile_19__2_,
         regBoiz_regfile_19__1_, regBoiz_regfile_19__0_,
         regBoiz_regfile_18__31_, regBoiz_regfile_18__30_,
         regBoiz_regfile_18__29_, regBoiz_regfile_18__28_,
         regBoiz_regfile_18__27_, regBoiz_regfile_18__26_,
         regBoiz_regfile_18__25_, regBoiz_regfile_18__24_,
         regBoiz_regfile_18__23_, regBoiz_regfile_18__22_,
         regBoiz_regfile_18__21_, regBoiz_regfile_18__20_,
         regBoiz_regfile_18__19_, regBoiz_regfile_18__18_,
         regBoiz_regfile_18__17_, regBoiz_regfile_18__16_,
         regBoiz_regfile_18__15_, regBoiz_regfile_18__14_,
         regBoiz_regfile_18__13_, regBoiz_regfile_18__12_,
         regBoiz_regfile_18__11_, regBoiz_regfile_18__10_,
         regBoiz_regfile_18__9_, regBoiz_regfile_18__8_,
         regBoiz_regfile_18__7_, regBoiz_regfile_18__6_,
         regBoiz_regfile_18__5_, regBoiz_regfile_18__4_,
         regBoiz_regfile_18__3_, regBoiz_regfile_18__2_,
         regBoiz_regfile_18__1_, regBoiz_regfile_18__0_,
         regBoiz_regfile_17__31_, regBoiz_regfile_17__30_,
         regBoiz_regfile_17__29_, regBoiz_regfile_17__28_,
         regBoiz_regfile_17__27_, regBoiz_regfile_17__26_,
         regBoiz_regfile_17__25_, regBoiz_regfile_17__24_,
         regBoiz_regfile_17__23_, regBoiz_regfile_17__22_,
         regBoiz_regfile_17__21_, regBoiz_regfile_17__20_,
         regBoiz_regfile_17__19_, regBoiz_regfile_17__18_,
         regBoiz_regfile_17__17_, regBoiz_regfile_17__16_,
         regBoiz_regfile_17__15_, regBoiz_regfile_17__14_,
         regBoiz_regfile_17__13_, regBoiz_regfile_17__12_,
         regBoiz_regfile_17__11_, regBoiz_regfile_17__10_,
         regBoiz_regfile_17__9_, regBoiz_regfile_17__8_,
         regBoiz_regfile_17__7_, regBoiz_regfile_17__6_,
         regBoiz_regfile_17__5_, regBoiz_regfile_17__4_,
         regBoiz_regfile_17__3_, regBoiz_regfile_17__2_,
         regBoiz_regfile_17__1_, regBoiz_regfile_17__0_,
         regBoiz_regfile_16__31_, regBoiz_regfile_16__30_,
         regBoiz_regfile_16__29_, regBoiz_regfile_16__28_,
         regBoiz_regfile_16__27_, regBoiz_regfile_16__26_,
         regBoiz_regfile_16__25_, regBoiz_regfile_16__24_,
         regBoiz_regfile_16__23_, regBoiz_regfile_16__22_,
         regBoiz_regfile_16__21_, regBoiz_regfile_16__20_,
         regBoiz_regfile_16__19_, regBoiz_regfile_16__18_,
         regBoiz_regfile_16__17_, regBoiz_regfile_16__16_,
         regBoiz_regfile_16__15_, regBoiz_regfile_16__14_,
         regBoiz_regfile_16__13_, regBoiz_regfile_16__12_,
         regBoiz_regfile_16__11_, regBoiz_regfile_16__10_,
         regBoiz_regfile_16__9_, regBoiz_regfile_16__8_,
         regBoiz_regfile_16__7_, regBoiz_regfile_16__6_,
         regBoiz_regfile_16__5_, regBoiz_regfile_16__4_,
         regBoiz_regfile_16__3_, regBoiz_regfile_16__2_,
         regBoiz_regfile_16__1_, regBoiz_regfile_16__0_,
         regBoiz_regfile_15__31_, regBoiz_regfile_15__30_,
         regBoiz_regfile_15__29_, regBoiz_regfile_15__28_,
         regBoiz_regfile_15__27_, regBoiz_regfile_15__26_,
         regBoiz_regfile_15__25_, regBoiz_regfile_15__24_,
         regBoiz_regfile_15__23_, regBoiz_regfile_15__22_,
         regBoiz_regfile_15__21_, regBoiz_regfile_15__20_,
         regBoiz_regfile_15__19_, regBoiz_regfile_15__18_,
         regBoiz_regfile_15__17_, regBoiz_regfile_15__16_,
         regBoiz_regfile_15__15_, regBoiz_regfile_15__14_,
         regBoiz_regfile_15__13_, regBoiz_regfile_15__12_,
         regBoiz_regfile_15__11_, regBoiz_regfile_15__10_,
         regBoiz_regfile_15__9_, regBoiz_regfile_15__8_,
         regBoiz_regfile_15__7_, regBoiz_regfile_15__6_,
         regBoiz_regfile_15__5_, regBoiz_regfile_15__4_,
         regBoiz_regfile_15__3_, regBoiz_regfile_15__2_,
         regBoiz_regfile_15__1_, regBoiz_regfile_15__0_,
         regBoiz_regfile_14__31_, regBoiz_regfile_14__30_,
         regBoiz_regfile_14__29_, regBoiz_regfile_14__28_,
         regBoiz_regfile_14__27_, regBoiz_regfile_14__26_,
         regBoiz_regfile_14__25_, regBoiz_regfile_14__24_,
         regBoiz_regfile_14__23_, regBoiz_regfile_14__22_,
         regBoiz_regfile_14__21_, regBoiz_regfile_14__20_,
         regBoiz_regfile_14__19_, regBoiz_regfile_14__18_,
         regBoiz_regfile_14__17_, regBoiz_regfile_14__16_,
         regBoiz_regfile_14__15_, regBoiz_regfile_14__14_,
         regBoiz_regfile_14__13_, regBoiz_regfile_14__12_,
         regBoiz_regfile_14__11_, regBoiz_regfile_14__10_,
         regBoiz_regfile_14__9_, regBoiz_regfile_14__8_,
         regBoiz_regfile_14__7_, regBoiz_regfile_14__6_,
         regBoiz_regfile_14__5_, regBoiz_regfile_14__4_,
         regBoiz_regfile_14__3_, regBoiz_regfile_14__2_,
         regBoiz_regfile_14__1_, regBoiz_regfile_14__0_,
         regBoiz_regfile_13__31_, regBoiz_regfile_13__30_,
         regBoiz_regfile_13__29_, regBoiz_regfile_13__28_,
         regBoiz_regfile_13__27_, regBoiz_regfile_13__26_,
         regBoiz_regfile_13__25_, regBoiz_regfile_13__24_,
         regBoiz_regfile_13__23_, regBoiz_regfile_13__22_,
         regBoiz_regfile_13__21_, regBoiz_regfile_13__20_,
         regBoiz_regfile_13__19_, regBoiz_regfile_13__18_,
         regBoiz_regfile_13__17_, regBoiz_regfile_13__16_,
         regBoiz_regfile_13__15_, regBoiz_regfile_13__14_,
         regBoiz_regfile_13__13_, regBoiz_regfile_13__12_,
         regBoiz_regfile_13__11_, regBoiz_regfile_13__10_,
         regBoiz_regfile_13__9_, regBoiz_regfile_13__8_,
         regBoiz_regfile_13__7_, regBoiz_regfile_13__6_,
         regBoiz_regfile_13__5_, regBoiz_regfile_13__4_,
         regBoiz_regfile_13__3_, regBoiz_regfile_13__2_,
         regBoiz_regfile_13__1_, regBoiz_regfile_13__0_,
         regBoiz_regfile_12__31_, regBoiz_regfile_12__30_,
         regBoiz_regfile_12__29_, regBoiz_regfile_12__28_,
         regBoiz_regfile_12__27_, regBoiz_regfile_12__26_,
         regBoiz_regfile_12__25_, regBoiz_regfile_12__24_,
         regBoiz_regfile_12__23_, regBoiz_regfile_12__22_,
         regBoiz_regfile_12__21_, regBoiz_regfile_12__20_,
         regBoiz_regfile_12__19_, regBoiz_regfile_12__18_,
         regBoiz_regfile_12__17_, regBoiz_regfile_12__16_,
         regBoiz_regfile_12__15_, regBoiz_regfile_12__14_,
         regBoiz_regfile_12__13_, regBoiz_regfile_12__12_,
         regBoiz_regfile_12__11_, regBoiz_regfile_12__10_,
         regBoiz_regfile_12__9_, regBoiz_regfile_12__8_,
         regBoiz_regfile_12__7_, regBoiz_regfile_12__6_,
         regBoiz_regfile_12__5_, regBoiz_regfile_12__4_,
         regBoiz_regfile_12__3_, regBoiz_regfile_12__2_,
         regBoiz_regfile_12__1_, regBoiz_regfile_12__0_,
         regBoiz_regfile_11__31_, regBoiz_regfile_11__30_,
         regBoiz_regfile_11__29_, regBoiz_regfile_11__28_,
         regBoiz_regfile_11__27_, regBoiz_regfile_11__26_,
         regBoiz_regfile_11__25_, regBoiz_regfile_11__24_,
         regBoiz_regfile_11__23_, regBoiz_regfile_11__22_,
         regBoiz_regfile_11__21_, regBoiz_regfile_11__20_,
         regBoiz_regfile_11__19_, regBoiz_regfile_11__18_,
         regBoiz_regfile_11__17_, regBoiz_regfile_11__16_,
         regBoiz_regfile_11__15_, regBoiz_regfile_11__14_,
         regBoiz_regfile_11__13_, regBoiz_regfile_11__12_,
         regBoiz_regfile_11__11_, regBoiz_regfile_11__10_,
         regBoiz_regfile_11__9_, regBoiz_regfile_11__8_,
         regBoiz_regfile_11__7_, regBoiz_regfile_11__6_,
         regBoiz_regfile_11__5_, regBoiz_regfile_11__4_,
         regBoiz_regfile_11__3_, regBoiz_regfile_11__2_,
         regBoiz_regfile_11__1_, regBoiz_regfile_11__0_,
         regBoiz_regfile_10__31_, regBoiz_regfile_10__30_,
         regBoiz_regfile_10__29_, regBoiz_regfile_10__28_,
         regBoiz_regfile_10__27_, regBoiz_regfile_10__26_,
         regBoiz_regfile_10__25_, regBoiz_regfile_10__24_,
         regBoiz_regfile_10__23_, regBoiz_regfile_10__22_,
         regBoiz_regfile_10__21_, regBoiz_regfile_10__20_,
         regBoiz_regfile_10__19_, regBoiz_regfile_10__18_,
         regBoiz_regfile_10__17_, regBoiz_regfile_10__16_,
         regBoiz_regfile_10__15_, regBoiz_regfile_10__14_,
         regBoiz_regfile_10__13_, regBoiz_regfile_10__12_,
         regBoiz_regfile_10__11_, regBoiz_regfile_10__10_,
         regBoiz_regfile_10__9_, regBoiz_regfile_10__8_,
         regBoiz_regfile_10__7_, regBoiz_regfile_10__6_,
         regBoiz_regfile_10__5_, regBoiz_regfile_10__4_,
         regBoiz_regfile_10__3_, regBoiz_regfile_10__2_,
         regBoiz_regfile_10__1_, regBoiz_regfile_10__0_,
         regBoiz_regfile_9__31_, regBoiz_regfile_9__30_,
         regBoiz_regfile_9__29_, regBoiz_regfile_9__28_,
         regBoiz_regfile_9__27_, regBoiz_regfile_9__26_,
         regBoiz_regfile_9__25_, regBoiz_regfile_9__24_,
         regBoiz_regfile_9__23_, regBoiz_regfile_9__22_,
         regBoiz_regfile_9__21_, regBoiz_regfile_9__20_,
         regBoiz_regfile_9__19_, regBoiz_regfile_9__18_,
         regBoiz_regfile_9__17_, regBoiz_regfile_9__16_,
         regBoiz_regfile_9__15_, regBoiz_regfile_9__14_,
         regBoiz_regfile_9__13_, regBoiz_regfile_9__12_,
         regBoiz_regfile_9__11_, regBoiz_regfile_9__10_, regBoiz_regfile_9__9_,
         regBoiz_regfile_9__8_, regBoiz_regfile_9__7_, regBoiz_regfile_9__6_,
         regBoiz_regfile_9__5_, regBoiz_regfile_9__4_, regBoiz_regfile_9__3_,
         regBoiz_regfile_9__2_, regBoiz_regfile_9__1_, regBoiz_regfile_9__0_,
         regBoiz_regfile_8__31_, regBoiz_regfile_8__30_,
         regBoiz_regfile_8__29_, regBoiz_regfile_8__28_,
         regBoiz_regfile_8__27_, regBoiz_regfile_8__26_,
         regBoiz_regfile_8__25_, regBoiz_regfile_8__24_,
         regBoiz_regfile_8__23_, regBoiz_regfile_8__22_,
         regBoiz_regfile_8__21_, regBoiz_regfile_8__20_,
         regBoiz_regfile_8__19_, regBoiz_regfile_8__18_,
         regBoiz_regfile_8__17_, regBoiz_regfile_8__16_,
         regBoiz_regfile_8__15_, regBoiz_regfile_8__14_,
         regBoiz_regfile_8__13_, regBoiz_regfile_8__12_,
         regBoiz_regfile_8__11_, regBoiz_regfile_8__10_, regBoiz_regfile_8__9_,
         regBoiz_regfile_8__8_, regBoiz_regfile_8__7_, regBoiz_regfile_8__6_,
         regBoiz_regfile_8__5_, regBoiz_regfile_8__4_, regBoiz_regfile_8__3_,
         regBoiz_regfile_8__2_, regBoiz_regfile_8__1_, regBoiz_regfile_8__0_,
         regBoiz_regfile_7__31_, regBoiz_regfile_7__30_,
         regBoiz_regfile_7__29_, regBoiz_regfile_7__28_,
         regBoiz_regfile_7__27_, regBoiz_regfile_7__26_,
         regBoiz_regfile_7__25_, regBoiz_regfile_7__24_,
         regBoiz_regfile_7__23_, regBoiz_regfile_7__22_,
         regBoiz_regfile_7__21_, regBoiz_regfile_7__20_,
         regBoiz_regfile_7__19_, regBoiz_regfile_7__18_,
         regBoiz_regfile_7__17_, regBoiz_regfile_7__16_,
         regBoiz_regfile_7__15_, regBoiz_regfile_7__14_,
         regBoiz_regfile_7__13_, regBoiz_regfile_7__12_,
         regBoiz_regfile_7__11_, regBoiz_regfile_7__10_, regBoiz_regfile_7__9_,
         regBoiz_regfile_7__8_, regBoiz_regfile_7__7_, regBoiz_regfile_7__6_,
         regBoiz_regfile_7__5_, regBoiz_regfile_7__4_, regBoiz_regfile_7__3_,
         regBoiz_regfile_7__2_, regBoiz_regfile_7__1_, regBoiz_regfile_7__0_,
         regBoiz_regfile_6__31_, regBoiz_regfile_6__30_,
         regBoiz_regfile_6__29_, regBoiz_regfile_6__28_,
         regBoiz_regfile_6__27_, regBoiz_regfile_6__26_,
         regBoiz_regfile_6__25_, regBoiz_regfile_6__24_,
         regBoiz_regfile_6__23_, regBoiz_regfile_6__22_,
         regBoiz_regfile_6__21_, regBoiz_regfile_6__20_,
         regBoiz_regfile_6__19_, regBoiz_regfile_6__18_,
         regBoiz_regfile_6__17_, regBoiz_regfile_6__16_,
         regBoiz_regfile_6__15_, regBoiz_regfile_6__14_,
         regBoiz_regfile_6__13_, regBoiz_regfile_6__12_,
         regBoiz_regfile_6__11_, regBoiz_regfile_6__10_, regBoiz_regfile_6__9_,
         regBoiz_regfile_6__8_, regBoiz_regfile_6__7_, regBoiz_regfile_6__6_,
         regBoiz_regfile_6__5_, regBoiz_regfile_6__4_, regBoiz_regfile_6__3_,
         regBoiz_regfile_6__2_, regBoiz_regfile_6__1_, regBoiz_regfile_6__0_,
         regBoiz_regfile_5__31_, regBoiz_regfile_5__30_,
         regBoiz_regfile_5__29_, regBoiz_regfile_5__28_,
         regBoiz_regfile_5__27_, regBoiz_regfile_5__26_,
         regBoiz_regfile_5__25_, regBoiz_regfile_5__24_,
         regBoiz_regfile_5__23_, regBoiz_regfile_5__22_,
         regBoiz_regfile_5__21_, regBoiz_regfile_5__20_,
         regBoiz_regfile_5__19_, regBoiz_regfile_5__18_,
         regBoiz_regfile_5__17_, regBoiz_regfile_5__16_,
         regBoiz_regfile_5__15_, regBoiz_regfile_5__14_,
         regBoiz_regfile_5__13_, regBoiz_regfile_5__12_,
         regBoiz_regfile_5__11_, regBoiz_regfile_5__10_, regBoiz_regfile_5__9_,
         regBoiz_regfile_5__8_, regBoiz_regfile_5__7_, regBoiz_regfile_5__6_,
         regBoiz_regfile_5__5_, regBoiz_regfile_5__4_, regBoiz_regfile_5__3_,
         regBoiz_regfile_5__2_, regBoiz_regfile_5__1_, regBoiz_regfile_5__0_,
         regBoiz_regfile_4__31_, regBoiz_regfile_4__30_,
         regBoiz_regfile_4__29_, regBoiz_regfile_4__28_,
         regBoiz_regfile_4__27_, regBoiz_regfile_4__26_,
         regBoiz_regfile_4__25_, regBoiz_regfile_4__24_,
         regBoiz_regfile_4__23_, regBoiz_regfile_4__22_,
         regBoiz_regfile_4__21_, regBoiz_regfile_4__20_,
         regBoiz_regfile_4__19_, regBoiz_regfile_4__18_,
         regBoiz_regfile_4__17_, regBoiz_regfile_4__16_,
         regBoiz_regfile_4__15_, regBoiz_regfile_4__14_,
         regBoiz_regfile_4__13_, regBoiz_regfile_4__12_,
         regBoiz_regfile_4__11_, regBoiz_regfile_4__10_, regBoiz_regfile_4__9_,
         regBoiz_regfile_4__8_, regBoiz_regfile_4__7_, regBoiz_regfile_4__6_,
         regBoiz_regfile_4__5_, regBoiz_regfile_4__4_, regBoiz_regfile_4__3_,
         regBoiz_regfile_4__2_, regBoiz_regfile_4__1_, regBoiz_regfile_4__0_,
         regBoiz_regfile_3__31_, regBoiz_regfile_3__30_,
         regBoiz_regfile_3__29_, regBoiz_regfile_3__28_,
         regBoiz_regfile_3__27_, regBoiz_regfile_3__26_,
         regBoiz_regfile_3__25_, regBoiz_regfile_3__24_,
         regBoiz_regfile_3__23_, regBoiz_regfile_3__22_,
         regBoiz_regfile_3__21_, regBoiz_regfile_3__20_,
         regBoiz_regfile_3__19_, regBoiz_regfile_3__18_,
         regBoiz_regfile_3__17_, regBoiz_regfile_3__16_,
         regBoiz_regfile_3__15_, regBoiz_regfile_3__14_,
         regBoiz_regfile_3__13_, regBoiz_regfile_3__12_,
         regBoiz_regfile_3__11_, regBoiz_regfile_3__10_, regBoiz_regfile_3__9_,
         regBoiz_regfile_3__8_, regBoiz_regfile_3__7_, regBoiz_regfile_3__6_,
         regBoiz_regfile_3__5_, regBoiz_regfile_3__4_, regBoiz_regfile_3__3_,
         regBoiz_regfile_3__2_, regBoiz_regfile_3__1_, regBoiz_regfile_3__0_,
         regBoiz_regfile_2__31_, regBoiz_regfile_2__30_,
         regBoiz_regfile_2__29_, regBoiz_regfile_2__28_,
         regBoiz_regfile_2__27_, regBoiz_regfile_2__26_,
         regBoiz_regfile_2__25_, regBoiz_regfile_2__24_,
         regBoiz_regfile_2__23_, regBoiz_regfile_2__22_,
         regBoiz_regfile_2__21_, regBoiz_regfile_2__20_,
         regBoiz_regfile_2__19_, regBoiz_regfile_2__18_,
         regBoiz_regfile_2__17_, regBoiz_regfile_2__16_,
         regBoiz_regfile_2__15_, regBoiz_regfile_2__14_,
         regBoiz_regfile_2__13_, regBoiz_regfile_2__12_,
         regBoiz_regfile_2__11_, regBoiz_regfile_2__10_, regBoiz_regfile_2__9_,
         regBoiz_regfile_2__8_, regBoiz_regfile_2__7_, regBoiz_regfile_2__6_,
         regBoiz_regfile_2__5_, regBoiz_regfile_2__4_, regBoiz_regfile_2__3_,
         regBoiz_regfile_2__2_, regBoiz_regfile_2__1_, regBoiz_regfile_2__0_,
         regBoiz_regfile_1__31_, regBoiz_regfile_1__30_,
         regBoiz_regfile_1__29_, regBoiz_regfile_1__28_,
         regBoiz_regfile_1__27_, regBoiz_regfile_1__26_,
         regBoiz_regfile_1__25_, regBoiz_regfile_1__24_,
         regBoiz_regfile_1__23_, regBoiz_regfile_1__22_,
         regBoiz_regfile_1__21_, regBoiz_regfile_1__20_,
         regBoiz_regfile_1__19_, regBoiz_regfile_1__18_,
         regBoiz_regfile_1__17_, regBoiz_regfile_1__16_,
         regBoiz_regfile_1__15_, regBoiz_regfile_1__14_,
         regBoiz_regfile_1__13_, regBoiz_regfile_1__12_,
         regBoiz_regfile_1__11_, regBoiz_regfile_1__10_, regBoiz_regfile_1__9_,
         regBoiz_regfile_1__8_, regBoiz_regfile_1__7_, regBoiz_regfile_1__6_,
         regBoiz_regfile_1__5_, regBoiz_regfile_1__4_, regBoiz_regfile_1__3_,
         regBoiz_regfile_1__2_, regBoiz_regfile_1__1_, regBoiz_regfile_1__0_,
         regBoiz_regfile_0__31_, regBoiz_regfile_0__30_,
         regBoiz_regfile_0__29_, regBoiz_regfile_0__28_,
         regBoiz_regfile_0__27_, regBoiz_regfile_0__26_,
         regBoiz_regfile_0__25_, regBoiz_regfile_0__24_,
         regBoiz_regfile_0__23_, regBoiz_regfile_0__22_,
         regBoiz_regfile_0__21_, regBoiz_regfile_0__20_,
         regBoiz_regfile_0__19_, regBoiz_regfile_0__18_,
         regBoiz_regfile_0__17_, regBoiz_regfile_0__16_,
         regBoiz_regfile_0__15_, regBoiz_regfile_0__14_,
         regBoiz_regfile_0__13_, regBoiz_regfile_0__12_,
         regBoiz_regfile_0__11_, regBoiz_regfile_0__10_, regBoiz_regfile_0__9_,
         regBoiz_regfile_0__8_, regBoiz_regfile_0__7_, regBoiz_regfile_0__6_,
         regBoiz_regfile_0__5_, regBoiz_regfile_0__4_, regBoiz_regfile_0__3_,
         regBoiz_regfile_0__2_, regBoiz_regfile_0__1_, regBoiz_regfile_0__0_,
         regBoiz_N18, regBoiz_N17, regBoiz_N16, regBoiz_N15, regBoiz_N12,
         aluBoi_condOut_0_, aluBoi_imm32w_0_, aluBoi_imm32w_1_,
         aluBoi_imm32w_2_, aluBoi_imm32w_3_, aluBoi_imm32w_4_,
         aluBoi_imm32w_5_, aluBoi_imm32w_6_, aluBoi_imm32w_7_,
         aluBoi_imm32w_8_, aluBoi_imm32w_9_, aluBoi_imm32w_10_,
         aluBoi_imm32w_11_, aluBoi_imm32w_12_, aluBoi_imm32w_13_,
         aluBoi_imm32w_14_, aluBoi_imm32w_15_, aluBoi_condBoi_N25,
         aluBoi_condBoi_N24, aluBoi_multBoi_N73, aluBoi_multBoi_N72,
         aluBoi_multBoi_N71, aluBoi_multBoi_N70, aluBoi_multBoi_N69,
         aluBoi_multBoi_N68, aluBoi_multBoi_N67, aluBoi_multBoi_N66,
         aluBoi_multBoi_N65, aluBoi_multBoi_N64, aluBoi_multBoi_N63,
         aluBoi_multBoi_N62, aluBoi_multBoi_N61, aluBoi_multBoi_N60,
         aluBoi_multBoi_N59, aluBoi_multBoi_N58, aluBoi_multBoi_N57,
         aluBoi_multBoi_N56, aluBoi_multBoi_N55, aluBoi_multBoi_N54,
         aluBoi_multBoi_N52, aluBoi_multBoi_N51, aluBoi_multBoi_N50,
         aluBoi_multBoi_N49, aluBoi_multBoi_N48, aluBoi_multBoi_N47,
         aluBoi_multBoi_N46, aluBoi_multBoi_N45, aluBoi_multBoi_N44,
         aluBoi_multBoi_N43, aluBoi_multBoi_N42, aluBoi_multBoi_N41,
         aluBoi_multBoi_N40, aluBoi_multBoi_N38, aluBoi_multBoi_N37,
         aluBoi_multBoi_N36, aluBoi_multBoi_N35, aluBoi_multBoi_N34,
         aluBoi_multBoi_N6, aluBoi_multBoi_count_0_, aluBoi_multBoi_count_1_,
         aluBoi_multBoi_count_2_, aluBoi_multBoi_runProd_0_, n34, n36, n38,
         n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62, n64, n66,
         n68, n70, n72, n74, n76, n78, n80, n82, n84, n86, n88, n90, n92, n94,
         n96, n98, n99, n100, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n607, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1145, n1146, n1147, n1149,
         n1151, n1153, n1157, n1158, n1162, n1165, n1168, n1171, n1174, n1177,
         n1180, n1183, n1186, n1189, n1192, n1195, n1198, n1201, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1213, n1214, n1216, n1219, n1221,
         n1223, n1225, n1227, n1229, n1232, n1234, n1236, n1238, n2009, n2010,
         n2011, n2013, n2014, n2054, n2082, n2105, n2202, n2203, n2204, n2840,
         n2841, n2842, n2844, n2847, n2983, n2984, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n3083, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3391, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4655, n4656, n4657, n4658, n4660, n4661, n4662,
         n4663, n4665, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4723, n4726, n4729, n4730, n4733, n4734, n4736, n4738,
         n4739, n4741, n4743, n4745, n4746, n4748, n4750, n4752, n4753, n4755,
         n4757, n4759, n4761, n4763, n4765, n4767, n4769, n4771, n4773, n4775,
         n4777, n4779, n4781, n4782, n4783, n4784, n4786, n4787, n4788, n4789,
         n4790, n4791, n4794, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4808, n4809, n4810, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4837, n4841, n4873, n4874,
         n4876, net129670, net327826, net328053, net329432, net334218,
         net345751, net358577, net358591, net358604, net358618, net359418,
         net359439, net359447, net359448, net359449, net359450, net359451,
         net359459, net359462, net359465, net359469, net359470, net359472,
         net359473, net359475, net359481, net359486, net359487, net359495,
         net359497, net359501, net359507, net359512, net359513, net359515,
         net359520, net359521, net359524, net359531, net359532, net359533,
         net359535, net359537, net359540, net359550, net359552, net359553,
         net359555, net359557, net359574, net359577, net359601, net359603,
         net359648, net359650, net359651, net359673, net359675, net359676,
         net359678, net359680, net359681, net359682, net359752, net359756,
         net359761, net359762, net359765, net359766, net359767, net359770,
         net359771, net359782, net359785, net359788, net359792, net359809,
         net359876, net359877, net359899, net359904, net359905, net359911,
         net359914, net359915, net359916, net359918, net359919, net359923,
         net359942, net359986, net360002, net360011, net360017, net360033,
         net360197, net360198, net360205, net360206, net360235, net360253,
         net360254, net360259, net360261, net360262, net360265, net360266,
         net360273, net360278, net360279, net360285, net360297, net360299,
         net360360, net360403, net360445, net360474, net360490, net360497,
         net360513, net360539, net360550, net360583, net360604, net360605,
         net360606, net360607, net360611, net360617, net360619, net360620,
         net360628, net360631, net360632, net360636, net360639, net360651,
         net360713, net360723, net360821, net360904, net360914, net360915,
         net360927, net360996, net361001, net361002, net361007, net361008,
         net361009, net361013, net361015, net361018, net361019, net361020,
         net361021, net361022, net361027, net361028, net361030, net361031,
         net361032, net361033, net361053, net361056, net361057, net361073,
         net361076, net361077, net361083, net361088, net361090, net361260,
         net361261, net361275, net361276, net361278, net361289, net361290,
         net361291, net361292, net361293, net361295, net361296, net361299,
         net361302, net361306, net361307, net361308, net361309, net361312,
         net361318, net361319, net361320, net361321, net361326, net361327,
         net361342, net361354, net361356, net361357, net361358, net361361,
         net361372, net361386, net361390, net361391, net361394, net361396,
         net361398, net361400, net361401, net361404, net361416, net361417,
         net361437, net361443, net361491, net361509, net361512, net361523,
         net361524, net361536, net361537, net361541, net361543, net361545,
         net361546, net361547, net361548, net361629, net361630, net361631,
         net361670, net361709, net361713, net361714, net361740, net361746,
         net361748, net361749, net361756, net361801, net361802, net361808,
         net361809, net361814, net361825, net361827, net361828, net361829,
         net361830, net361833, net361835, net361838, net361885, net361886,
         net361889, net361890, net361891, net361893, net361899, net361900,
         net361902, net361903, net361906, net361907, net361911, net361913,
         net361949, net361984, net362016, net362026, net362028, net362047,
         net362048, net362049, net362050, net362052, net362053, net362061,
         net362062, net362091, net362092, net362094, net362095, net362096,
         net362097, net362105, net362107, net362108, net362109, net362110,
         net362117, net362122, net362124, net362125, net362126, net362127,
         net362131, net362134, net362141, net362142, net362146, net362149,
         net362152, net362153, net362156, net362157, net362158, net362159,
         net362161, net362172, net362175, net362177, net362178, net362179,
         net362194, net362196, net362211, net362216, net362218, net362223,
         net362224, net362229, net362230, net362231, net362233, net362238,
         net362239, net362240, net362246, net362251, net362253, net362255,
         net362256, net362257, net362262, net362265, net362269, net362270,
         net362281, net362287, net362297, net362311, net362312, net362314,
         net362317, net362318, net362322, net362327, net362330, net362337,
         net362341, net362342, net362361, net362362, net362387, net362485,
         net363046, net363047, net363049, net363057, net364246, net364764,
         net364779, net364803, net364870, net364871, net364874, net364875,
         net364882, net364898, net364899, net364904, net364905, net364906,
         net364941, net364968, net364970, net364971, net365030, net365031,
         net365032, net365033, net365093, net365099, net365100, net365106,
         net365284, net365293, net365335, net365336, net365399, net365830,
         net366184, net366907, net366905, net366901, net366899, net366887,
         net366885, net366953, net366951, net366949, net366947, net366945,
         net366939, net366937, net366935, net366933, net366927, net366925,
         net366923, net366921, net366919, net367009, net367007, net367005,
         net367003, net367001, net366999, net366997, net366995, net366991,
         net366987, net366985, net366981, net366979, net366977, net366973,
         net366971, net366969, net366967, net366965, net367045, net367043,
         net367041, net367039, net367035, net367031, net367029, net367027,
         net367025, net367023, net367019, net367221, net367217, net367215,
         net367231, net367597, net367595, net367593, net367631, net368069,
         net368183, net368181, net368179, net368187, net368185, net368201,
         net368195, net368205, net368203, net368215, net368213, net368211,
         net368209, net368217, net368225, net368223, net368221, net368436,
         net368447, net368446, net368445, net368444, net368442, net368462,
         net368461, net368467, net368498, net368502, net368501, net368519,
         net368548, net368572, net368571, net368584, net368583, net368676,
         net368681, net368713, net368712, net368782, net368781, net368787,
         net368800, net368862, net368903, net368927, net368926, net369096,
         net369137, net369166, net369165, net369164, net369163, net369162,
         net369161, net369160, net369158, net369157, net369156, net369155,
         net369154, net369149, net369148, net369147, net369145, net369144,
         net369143, net369142, net369140, net369139, net369138, net369197,
         net369210, net369208, net369206, net369204, net369202, net369200,
         net369216, net369214, net369212, net369224, net369222, net369220,
         net369218, net369232, net369230, net369228, net369226, net369240,
         net369236, net369234, net369248, net369246, net369244, net369242,
         net369287, net369286, net369316, net375279, net375310, net375309,
         net375336, net375393, net375435, net375434, net375506, net375510,
         net375528, net375527, net375526, net375525, net375547, net375614,
         net375618, net375642, net375650, net375713, net375718, net375717,
         net375721, net375727, net375738, net375769, net375768, net375794,
         net375793, net375867, net375876, net375929, net375948, net375980,
         net375993, net376063, net376077, net376076, net376121, net376223,
         net376222, net376322, net376321, net376331, net376330, net376374,
         net376387, net376417, net376541, net376574, net376579, net376602,
         net376642, net376691, net376785, net376800, net376879, net376877,
         net376916, net376914, net376961, net376960, net377071, net377133,
         net377166, net377338, net377337, net377355, net377373, net377444,
         net377443, net377452, net377454, net377453, net377462, net377464,
         net377501, net377513, net377531, net377575, net377576, net377607,
         net377611, net377689, net377695, net377700, net377791, net377800,
         net377817, net377909, net377937, net377947, net377979, net378013,
         net378052, net378060, net378128, net378138, net378137, net378220,
         net378318, net378321, net378368, net378405, net378422, net378488,
         net378491, net378494, net377481, net361410, net377900, net359772,
         net359679, net359474, net368518, net368435, net361080, net359754,
         net100474, net362139, net362138, net362063, net362051, net361411,
         net361081, net360015, net360014, net360003, net359504, net378432,
         net377530, net362113, net362112, net361834, net361029, net361025,
         net361023, net360926, net360618, net361263, net361262, net360626,
         net377081, net377080, net368497, net362232, net351631, net377375,
         net361335, net361325, net361324, net361322, net361270, net362140,
         net377660, net377502, net361277, net361271, net361268, net361266,
         net361265, net361264, net359784, net359783, net359554, net378103,
         net362323, net362321, net362136, net362135, net362130, net362121,
         net362120, net362116, net362114, net360004, net359492, net377550,
         net361409, net361279, net361274, net361273, net361272, net361079,
         net360005, net359471, net368547, net368466, net362268, net362266,
         net362264, net362237, net359966, net377784, net377602, net368481,
         net359652, net359499, net359494, net359493, net359490, net359489,
         net359488, net100619, net377824, net375910, net377109, net366911,
         net365095, net365087, net362286, net368775, net367013, net367011,
         net366993, net366989, net365091, net365090, net365089, net365088,
         net378336, net369285, net368191, net361511, net361510, net361380,
         net359750, net368440, net368439, net368786, net368770, net378420,
         net377383, net376826, net376139, net362166, net361832, net361831,
         net361535, net361532, net377342, net360288, net360287, net360283,
         net360282, net360008, net360007, net360006, net360635, net360634,
         net360284, net359913, net376582, net376581, net361006, net361000,
         net360919, net360633, net360629, net360625, net360623, net360621,
         net360609, net360608, net375305, net375304, net361539, net361530,
         net361529, net361526, net361433, net361387, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5011,
         n5012, n5014, n5015, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5750, n5751, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5765, n5766, n5767, n5768, n5769, n5770, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5982, n5983, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6266, n6267, n6268, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6279, n6280, n6281,
         n6282, n6283, n6284, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6374, n6375, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6395, n6396, n6399, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13538, n13539, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, aluBoi_aluBoi_shft_SRA_sra_25_n185,
         aluBoi_aluBoi_shft_SRA_sra_25_n184,
         aluBoi_aluBoi_shft_SRA_sra_25_n183,
         aluBoi_aluBoi_shft_SRA_sra_25_n182,
         aluBoi_aluBoi_shft_SRA_sra_25_n181,
         aluBoi_aluBoi_shft_SRA_sra_25_n180,
         aluBoi_aluBoi_shft_SRA_sra_25_n179,
         aluBoi_aluBoi_shft_SRA_sra_25_n178,
         aluBoi_aluBoi_shft_SRA_sra_25_n177,
         aluBoi_aluBoi_shft_SRA_sra_25_n176,
         aluBoi_aluBoi_shft_SRA_sra_25_n175,
         aluBoi_aluBoi_shft_SRA_sra_25_n174,
         aluBoi_aluBoi_shft_SRA_sra_25_n173,
         aluBoi_aluBoi_shft_SRA_sra_25_n172,
         aluBoi_aluBoi_shft_SRA_sra_25_n171,
         aluBoi_aluBoi_shft_SRA_sra_25_n170,
         aluBoi_aluBoi_shft_SRA_sra_25_n169,
         aluBoi_aluBoi_shft_SRA_sra_25_n168,
         aluBoi_aluBoi_shft_SRA_sra_25_n167,
         aluBoi_aluBoi_shft_SRA_sra_25_n166,
         aluBoi_aluBoi_shft_SRA_sra_25_n165,
         aluBoi_aluBoi_shft_SRA_sra_25_n164,
         aluBoi_aluBoi_shft_SRA_sra_25_n163,
         aluBoi_aluBoi_shft_SRA_sra_25_n162,
         aluBoi_aluBoi_shft_SRA_sra_25_n161,
         aluBoi_aluBoi_shft_SRA_sra_25_n160,
         aluBoi_aluBoi_shft_SRA_sra_25_n159,
         aluBoi_aluBoi_shft_SRA_sra_25_n158,
         aluBoi_aluBoi_shft_SRA_sra_25_n157,
         aluBoi_aluBoi_shft_SRA_sra_25_n156,
         aluBoi_aluBoi_shft_SRA_sra_25_n155,
         aluBoi_aluBoi_shft_SRA_sra_25_n154,
         aluBoi_aluBoi_shft_SRA_sra_25_n153,
         aluBoi_aluBoi_shft_SRA_sra_25_n152,
         aluBoi_aluBoi_shft_SRA_sra_25_n151,
         aluBoi_aluBoi_shft_SRA_sra_25_n150,
         aluBoi_aluBoi_shft_SRA_sra_25_n149,
         aluBoi_aluBoi_shft_SRA_sra_25_n148,
         aluBoi_aluBoi_shft_SRA_sra_25_n147,
         aluBoi_aluBoi_shft_SRA_sra_25_n146,
         aluBoi_aluBoi_shft_SRA_sra_25_n145,
         aluBoi_aluBoi_shft_SRA_sra_25_n144,
         aluBoi_aluBoi_shft_SRA_sra_25_n143,
         aluBoi_aluBoi_shft_SRA_sra_25_n142,
         aluBoi_aluBoi_shft_SRA_sra_25_n141,
         aluBoi_aluBoi_shft_SRA_sra_25_n140,
         aluBoi_aluBoi_shft_SRA_sra_25_n139,
         aluBoi_aluBoi_shft_SRA_sra_25_n138,
         aluBoi_aluBoi_shft_SRA_sra_25_n137,
         aluBoi_aluBoi_shft_SRA_sra_25_n136,
         aluBoi_aluBoi_shft_SRA_sra_25_n135,
         aluBoi_aluBoi_shft_SRA_sra_25_n134,
         aluBoi_aluBoi_shft_SRA_sra_25_n133,
         aluBoi_aluBoi_shft_SRA_sra_25_n132,
         aluBoi_aluBoi_shft_SRA_sra_25_n131,
         aluBoi_aluBoi_shft_SRA_sra_25_n130,
         aluBoi_aluBoi_shft_SRA_sra_25_n129,
         aluBoi_aluBoi_shft_SRA_sra_25_n128,
         aluBoi_aluBoi_shft_SRA_sra_25_n127,
         aluBoi_aluBoi_shft_SRA_sra_25_n126,
         aluBoi_aluBoi_shft_SRA_sra_25_n125,
         aluBoi_aluBoi_shft_SRA_sra_25_n124,
         aluBoi_aluBoi_shft_SRA_sra_25_n123,
         aluBoi_aluBoi_shft_SRA_sra_25_n122,
         aluBoi_aluBoi_shft_SRA_sra_25_n121,
         aluBoi_aluBoi_shft_SRA_sra_25_n120,
         aluBoi_aluBoi_shft_SRA_sra_25_n119,
         aluBoi_aluBoi_shft_SRA_sra_25_n118,
         aluBoi_aluBoi_shft_SRA_sra_25_n117,
         aluBoi_aluBoi_shft_SRA_sra_25_n116,
         aluBoi_aluBoi_shft_SRA_sra_25_n115,
         aluBoi_aluBoi_shft_SRA_sra_25_n114,
         aluBoi_aluBoi_shft_SRA_sra_25_n113,
         aluBoi_aluBoi_shft_SRA_sra_25_n112,
         aluBoi_aluBoi_shft_SRA_sra_25_n111,
         aluBoi_aluBoi_shft_SRA_sra_25_n110,
         aluBoi_aluBoi_shft_SRA_sra_25_n109,
         aluBoi_aluBoi_shft_SRA_sra_25_n108,
         aluBoi_aluBoi_shft_SRA_sra_25_n107,
         aluBoi_aluBoi_shft_SRA_sra_25_n106,
         aluBoi_aluBoi_shft_SRA_sra_25_n105,
         aluBoi_aluBoi_shft_SRA_sra_25_n104,
         aluBoi_aluBoi_shft_SRA_sra_25_n103,
         aluBoi_aluBoi_shft_SRA_sra_25_n102,
         aluBoi_aluBoi_shft_SRA_sra_25_n101,
         aluBoi_aluBoi_shft_SRA_sra_25_n100, aluBoi_aluBoi_shft_SRA_sra_25_n99,
         aluBoi_aluBoi_shft_SRA_sra_25_n98, aluBoi_aluBoi_shft_SRA_sra_25_n97,
         aluBoi_aluBoi_shft_SRA_sra_25_n96, aluBoi_aluBoi_shft_SRA_sra_25_n95,
         aluBoi_aluBoi_shft_SRA_sra_25_n94, aluBoi_aluBoi_shft_SRA_sra_25_n93,
         aluBoi_aluBoi_shft_SRA_sra_25_n92, aluBoi_aluBoi_shft_SRA_sra_25_n91,
         aluBoi_aluBoi_shft_SRA_sra_25_n90, aluBoi_aluBoi_shft_SRA_sra_25_n89,
         aluBoi_aluBoi_shft_SRA_sra_25_n88, aluBoi_aluBoi_shft_SRA_sra_25_n87,
         aluBoi_aluBoi_shft_SRA_sra_25_n86, aluBoi_aluBoi_shft_SRA_sra_25_n85,
         aluBoi_aluBoi_shft_SRA_sra_25_n84, aluBoi_aluBoi_shft_SRA_sra_25_n83,
         aluBoi_aluBoi_shft_SRA_sra_25_n82, aluBoi_aluBoi_shft_SRA_sra_25_n81,
         aluBoi_aluBoi_shft_SRA_sra_25_n80, aluBoi_aluBoi_shft_SRA_sra_25_n79,
         aluBoi_aluBoi_shft_SRA_sra_25_n78, aluBoi_aluBoi_shft_SRA_sra_25_n77,
         aluBoi_aluBoi_shft_SRA_sra_25_n76, aluBoi_aluBoi_shft_SRA_sra_25_n75,
         aluBoi_aluBoi_shft_SRA_sra_25_n74, aluBoi_aluBoi_shft_SRA_sra_25_n73,
         aluBoi_aluBoi_shft_SRA_sra_25_n72, aluBoi_aluBoi_shft_SRA_sra_25_n71,
         aluBoi_aluBoi_shft_SRA_sra_25_n70, aluBoi_aluBoi_shft_SRA_sra_25_n69,
         aluBoi_aluBoi_shft_SRA_sra_25_n68, aluBoi_aluBoi_shft_SRA_sra_25_n67,
         aluBoi_aluBoi_shft_SRA_sra_25_n66, aluBoi_aluBoi_shft_SRA_sra_25_n65,
         aluBoi_aluBoi_shft_SRA_sra_25_n64, aluBoi_aluBoi_shft_SRA_sra_25_n63,
         aluBoi_aluBoi_shft_SRA_sra_25_n62, aluBoi_aluBoi_shft_SRA_sra_25_n61,
         aluBoi_aluBoi_shft_SRA_sra_25_n60, aluBoi_aluBoi_shft_SRA_sra_25_n59,
         aluBoi_aluBoi_shft_SRA_sra_25_n58, aluBoi_aluBoi_shft_SRA_sra_25_n57,
         aluBoi_aluBoi_shft_SRA_sra_25_n56, aluBoi_aluBoi_shft_SRA_sra_25_n55,
         aluBoi_aluBoi_shft_SRA_sra_25_n54, aluBoi_aluBoi_shft_SRA_sra_25_n53,
         aluBoi_aluBoi_shft_SRA_sra_25_n52, aluBoi_aluBoi_shft_SRA_sra_25_n51,
         aluBoi_aluBoi_shft_SRA_sra_25_n50, aluBoi_aluBoi_shft_SRA_sra_25_n49,
         aluBoi_aluBoi_shft_SRA_sra_25_n48, aluBoi_aluBoi_shft_SRA_sra_25_n47,
         aluBoi_aluBoi_shft_SRA_sra_25_n46, aluBoi_aluBoi_shft_SRA_sra_25_n45,
         aluBoi_aluBoi_shft_SRA_sra_25_n44, aluBoi_aluBoi_shft_SRA_sra_25_n43,
         aluBoi_aluBoi_shft_SRA_sra_25_n42, aluBoi_aluBoi_shft_SRA_sra_25_n41,
         aluBoi_aluBoi_shft_SRA_sra_25_n40, aluBoi_aluBoi_shft_SRA_sra_25_n39,
         aluBoi_aluBoi_shft_SRA_sra_25_n38, aluBoi_aluBoi_shft_SRA_sra_25_n37,
         aluBoi_aluBoi_shft_SRA_sra_25_n36, aluBoi_aluBoi_shft_SRA_sra_25_n35,
         aluBoi_aluBoi_shft_SRA_sra_25_n34, aluBoi_aluBoi_shft_SRA_sra_25_n33,
         aluBoi_aluBoi_shft_SRA_sra_25_n32, aluBoi_aluBoi_shft_SRA_sra_25_n31,
         aluBoi_aluBoi_shft_SRA_sra_25_n30, aluBoi_aluBoi_shft_SRA_sra_25_n29,
         aluBoi_aluBoi_shft_SRA_sra_25_n28, aluBoi_aluBoi_shft_SRA_sra_25_n27,
         aluBoi_aluBoi_shft_SRA_sra_25_n26, aluBoi_aluBoi_shft_SRA_sra_25_n25,
         aluBoi_aluBoi_shft_SRA_sra_25_n24, aluBoi_aluBoi_shft_SRA_sra_25_n23,
         aluBoi_aluBoi_shft_SRA_sra_25_n22, aluBoi_aluBoi_shft_SRA_sra_25_n21,
         aluBoi_aluBoi_shft_SRA_sra_25_n20, aluBoi_aluBoi_shft_SRA_sra_25_n19,
         aluBoi_aluBoi_shft_SRA_sra_25_n18, aluBoi_aluBoi_shft_SRA_sra_25_n17,
         aluBoi_aluBoi_shft_SRA_sra_25_n16, aluBoi_aluBoi_shft_SRA_sra_25_n15,
         aluBoi_aluBoi_shft_SRA_sra_25_n14, aluBoi_aluBoi_shft_SRA_sra_25_n13,
         aluBoi_aluBoi_shft_SRA_sra_25_n12, aluBoi_aluBoi_shft_SRA_sra_25_n11,
         aluBoi_aluBoi_shft_SRA_sra_25_n10, aluBoi_aluBoi_shft_SRA_sra_25_n9,
         aluBoi_aluBoi_shft_SRA_sra_25_n8, aluBoi_aluBoi_shft_SRA_sra_25_n7,
         aluBoi_aluBoi_shft_SRA_sra_25_n6, aluBoi_aluBoi_shft_SRA_sra_25_n5,
         aluBoi_aluBoi_shft_SRA_sra_25_n4, aluBoi_aluBoi_shft_SRA_sra_25_n3,
         aluBoi_aluBoi_shft_SRA_sra_25_n2, aluBoi_aluBoi_shft_SRA_sra_25_n1,
         aluBoi_aluBoi_shft_SRL_srl_16_n184,
         aluBoi_aluBoi_shft_SRL_srl_16_n183,
         aluBoi_aluBoi_shft_SRL_srl_16_n182,
         aluBoi_aluBoi_shft_SRL_srl_16_n181,
         aluBoi_aluBoi_shft_SRL_srl_16_n180,
         aluBoi_aluBoi_shft_SRL_srl_16_n179,
         aluBoi_aluBoi_shft_SRL_srl_16_n178,
         aluBoi_aluBoi_shft_SRL_srl_16_n177,
         aluBoi_aluBoi_shft_SRL_srl_16_n176,
         aluBoi_aluBoi_shft_SRL_srl_16_n175,
         aluBoi_aluBoi_shft_SRL_srl_16_n174,
         aluBoi_aluBoi_shft_SRL_srl_16_n173,
         aluBoi_aluBoi_shft_SRL_srl_16_n172,
         aluBoi_aluBoi_shft_SRL_srl_16_n171,
         aluBoi_aluBoi_shft_SRL_srl_16_n170,
         aluBoi_aluBoi_shft_SRL_srl_16_n169,
         aluBoi_aluBoi_shft_SRL_srl_16_n168,
         aluBoi_aluBoi_shft_SRL_srl_16_n167,
         aluBoi_aluBoi_shft_SRL_srl_16_n166,
         aluBoi_aluBoi_shft_SRL_srl_16_n165,
         aluBoi_aluBoi_shft_SRL_srl_16_n164,
         aluBoi_aluBoi_shft_SRL_srl_16_n163,
         aluBoi_aluBoi_shft_SRL_srl_16_n162,
         aluBoi_aluBoi_shft_SRL_srl_16_n161,
         aluBoi_aluBoi_shft_SRL_srl_16_n160,
         aluBoi_aluBoi_shft_SRL_srl_16_n159,
         aluBoi_aluBoi_shft_SRL_srl_16_n158,
         aluBoi_aluBoi_shft_SRL_srl_16_n157,
         aluBoi_aluBoi_shft_SRL_srl_16_n156,
         aluBoi_aluBoi_shft_SRL_srl_16_n155,
         aluBoi_aluBoi_shft_SRL_srl_16_n154,
         aluBoi_aluBoi_shft_SRL_srl_16_n153,
         aluBoi_aluBoi_shft_SRL_srl_16_n152,
         aluBoi_aluBoi_shft_SRL_srl_16_n151,
         aluBoi_aluBoi_shft_SRL_srl_16_n150,
         aluBoi_aluBoi_shft_SRL_srl_16_n149,
         aluBoi_aluBoi_shft_SRL_srl_16_n148,
         aluBoi_aluBoi_shft_SRL_srl_16_n147,
         aluBoi_aluBoi_shft_SRL_srl_16_n146,
         aluBoi_aluBoi_shft_SRL_srl_16_n145,
         aluBoi_aluBoi_shft_SRL_srl_16_n144,
         aluBoi_aluBoi_shft_SRL_srl_16_n143,
         aluBoi_aluBoi_shft_SRL_srl_16_n142,
         aluBoi_aluBoi_shft_SRL_srl_16_n141,
         aluBoi_aluBoi_shft_SRL_srl_16_n140,
         aluBoi_aluBoi_shft_SRL_srl_16_n139,
         aluBoi_aluBoi_shft_SRL_srl_16_n138,
         aluBoi_aluBoi_shft_SRL_srl_16_n137,
         aluBoi_aluBoi_shft_SRL_srl_16_n136,
         aluBoi_aluBoi_shft_SRL_srl_16_n135,
         aluBoi_aluBoi_shft_SRL_srl_16_n134,
         aluBoi_aluBoi_shft_SRL_srl_16_n133,
         aluBoi_aluBoi_shft_SRL_srl_16_n132,
         aluBoi_aluBoi_shft_SRL_srl_16_n131,
         aluBoi_aluBoi_shft_SRL_srl_16_n130,
         aluBoi_aluBoi_shft_SRL_srl_16_n129,
         aluBoi_aluBoi_shft_SRL_srl_16_n128,
         aluBoi_aluBoi_shft_SRL_srl_16_n127,
         aluBoi_aluBoi_shft_SRL_srl_16_n126,
         aluBoi_aluBoi_shft_SRL_srl_16_n125,
         aluBoi_aluBoi_shft_SRL_srl_16_n124,
         aluBoi_aluBoi_shft_SRL_srl_16_n123,
         aluBoi_aluBoi_shft_SRL_srl_16_n122,
         aluBoi_aluBoi_shft_SRL_srl_16_n121,
         aluBoi_aluBoi_shft_SRL_srl_16_n120,
         aluBoi_aluBoi_shft_SRL_srl_16_n119,
         aluBoi_aluBoi_shft_SRL_srl_16_n118,
         aluBoi_aluBoi_shft_SRL_srl_16_n117,
         aluBoi_aluBoi_shft_SRL_srl_16_n116,
         aluBoi_aluBoi_shft_SRL_srl_16_n115,
         aluBoi_aluBoi_shft_SRL_srl_16_n114,
         aluBoi_aluBoi_shft_SRL_srl_16_n113,
         aluBoi_aluBoi_shft_SRL_srl_16_n112,
         aluBoi_aluBoi_shft_SRL_srl_16_n111,
         aluBoi_aluBoi_shft_SRL_srl_16_n110,
         aluBoi_aluBoi_shft_SRL_srl_16_n109,
         aluBoi_aluBoi_shft_SRL_srl_16_n108,
         aluBoi_aluBoi_shft_SRL_srl_16_n107,
         aluBoi_aluBoi_shft_SRL_srl_16_n106,
         aluBoi_aluBoi_shft_SRL_srl_16_n105,
         aluBoi_aluBoi_shft_SRL_srl_16_n104,
         aluBoi_aluBoi_shft_SRL_srl_16_n103,
         aluBoi_aluBoi_shft_SRL_srl_16_n102,
         aluBoi_aluBoi_shft_SRL_srl_16_n101,
         aluBoi_aluBoi_shft_SRL_srl_16_n100, aluBoi_aluBoi_shft_SRL_srl_16_n99,
         aluBoi_aluBoi_shft_SRL_srl_16_n98, aluBoi_aluBoi_shft_SRL_srl_16_n97,
         aluBoi_aluBoi_shft_SRL_srl_16_n96, aluBoi_aluBoi_shft_SRL_srl_16_n95,
         aluBoi_aluBoi_shft_SRL_srl_16_n94, aluBoi_aluBoi_shft_SRL_srl_16_n93,
         aluBoi_aluBoi_shft_SRL_srl_16_n92, aluBoi_aluBoi_shft_SRL_srl_16_n91,
         aluBoi_aluBoi_shft_SRL_srl_16_n90, aluBoi_aluBoi_shft_SRL_srl_16_n89,
         aluBoi_aluBoi_shft_SRL_srl_16_n88, aluBoi_aluBoi_shft_SRL_srl_16_n87,
         aluBoi_aluBoi_shft_SRL_srl_16_n86, aluBoi_aluBoi_shft_SRL_srl_16_n85,
         aluBoi_aluBoi_shft_SRL_srl_16_n84, aluBoi_aluBoi_shft_SRL_srl_16_n83,
         aluBoi_aluBoi_shft_SRL_srl_16_n82, aluBoi_aluBoi_shft_SRL_srl_16_n81,
         aluBoi_aluBoi_shft_SRL_srl_16_n80, aluBoi_aluBoi_shft_SRL_srl_16_n79,
         aluBoi_aluBoi_shft_SRL_srl_16_n78, aluBoi_aluBoi_shft_SRL_srl_16_n77,
         aluBoi_aluBoi_shft_SRL_srl_16_n76, aluBoi_aluBoi_shft_SRL_srl_16_n75,
         aluBoi_aluBoi_shft_SRL_srl_16_n74, aluBoi_aluBoi_shft_SRL_srl_16_n73,
         aluBoi_aluBoi_shft_SRL_srl_16_n72, aluBoi_aluBoi_shft_SRL_srl_16_n71,
         aluBoi_aluBoi_shft_SRL_srl_16_n70, aluBoi_aluBoi_shft_SRL_srl_16_n69,
         aluBoi_aluBoi_shft_SRL_srl_16_n68, aluBoi_aluBoi_shft_SRL_srl_16_n67,
         aluBoi_aluBoi_shft_SRL_srl_16_n66, aluBoi_aluBoi_shft_SRL_srl_16_n65,
         aluBoi_aluBoi_shft_SRL_srl_16_n64, aluBoi_aluBoi_shft_SRL_srl_16_n63,
         aluBoi_aluBoi_shft_SRL_srl_16_n62, aluBoi_aluBoi_shft_SRL_srl_16_n61,
         aluBoi_aluBoi_shft_SRL_srl_16_n60, aluBoi_aluBoi_shft_SRL_srl_16_n59,
         aluBoi_aluBoi_shft_SRL_srl_16_n58, aluBoi_aluBoi_shft_SRL_srl_16_n57,
         aluBoi_aluBoi_shft_SRL_srl_16_n56, aluBoi_aluBoi_shft_SRL_srl_16_n55,
         aluBoi_aluBoi_shft_SRL_srl_16_n54, aluBoi_aluBoi_shft_SRL_srl_16_n53,
         aluBoi_aluBoi_shft_SRL_srl_16_n52, aluBoi_aluBoi_shft_SRL_srl_16_n51,
         aluBoi_aluBoi_shft_SRL_srl_16_n50, aluBoi_aluBoi_shft_SRL_srl_16_n49,
         aluBoi_aluBoi_shft_SRL_srl_16_n48, aluBoi_aluBoi_shft_SRL_srl_16_n47,
         aluBoi_aluBoi_shft_SRL_srl_16_n46, aluBoi_aluBoi_shft_SRL_srl_16_n45,
         aluBoi_aluBoi_shft_SRL_srl_16_n44, aluBoi_aluBoi_shft_SRL_srl_16_n43,
         aluBoi_aluBoi_shft_SRL_srl_16_n42, aluBoi_aluBoi_shft_SRL_srl_16_n41,
         aluBoi_aluBoi_shft_SRL_srl_16_n40, aluBoi_aluBoi_shft_SRL_srl_16_n39,
         aluBoi_aluBoi_shft_SRL_srl_16_n38, aluBoi_aluBoi_shft_SRL_srl_16_n37,
         aluBoi_aluBoi_shft_SRL_srl_16_n36, aluBoi_aluBoi_shft_SRL_srl_16_n35,
         aluBoi_aluBoi_shft_SRL_srl_16_n34, aluBoi_aluBoi_shft_SRL_srl_16_n33,
         aluBoi_aluBoi_shft_SRL_srl_16_n32, aluBoi_aluBoi_shft_SRL_srl_16_n31,
         aluBoi_aluBoi_shft_SRL_srl_16_n30, aluBoi_aluBoi_shft_SRL_srl_16_n28,
         aluBoi_aluBoi_shft_SRL_srl_16_n27, aluBoi_aluBoi_shft_SRL_srl_16_n26,
         aluBoi_aluBoi_shft_SRL_srl_16_n24, aluBoi_aluBoi_shft_SRL_srl_16_n22,
         aluBoi_aluBoi_shft_SRL_srl_16_n21, aluBoi_aluBoi_shft_SRL_srl_16_n20,
         aluBoi_aluBoi_shft_SRL_srl_16_n19, aluBoi_aluBoi_shft_SRL_srl_16_n18,
         aluBoi_aluBoi_shft_SRL_srl_16_n17, aluBoi_aluBoi_shft_SRL_srl_16_n16,
         aluBoi_aluBoi_shft_SRL_srl_16_n15, aluBoi_aluBoi_shft_SRL_srl_16_n14,
         aluBoi_aluBoi_shft_SRL_srl_16_n13, aluBoi_aluBoi_shft_SRL_srl_16_n12,
         aluBoi_aluBoi_shft_SRL_srl_16_n11, aluBoi_aluBoi_shft_SRL_srl_16_n10,
         aluBoi_aluBoi_shft_SRL_srl_16_n9, aluBoi_aluBoi_shft_SRL_srl_16_n8,
         aluBoi_aluBoi_shft_SRL_srl_16_n7, aluBoi_aluBoi_shft_SRL_srl_16_n6,
         aluBoi_aluBoi_shft_SRL_srl_16_n5, aluBoi_aluBoi_shft_SRL_srl_16_n4,
         aluBoi_aluBoi_shft_SRL_srl_16_n3, aluBoi_aluBoi_shft_SRL_srl_16_n2,
         aluBoi_aluBoi_shft_SRL_srl_16_n1, aluBoi_aluBoi_shft_SLL_sll_7_n40,
         aluBoi_aluBoi_shft_SLL_sll_7_n39, aluBoi_aluBoi_shft_SLL_sll_7_n38,
         aluBoi_aluBoi_shft_SLL_sll_7_n37, aluBoi_aluBoi_shft_SLL_sll_7_n36,
         aluBoi_aluBoi_shft_SLL_sll_7_n35, aluBoi_aluBoi_shft_SLL_sll_7_n34,
         aluBoi_aluBoi_shft_SLL_sll_7_n33, aluBoi_aluBoi_shft_SLL_sll_7_n32,
         aluBoi_aluBoi_shft_SLL_sll_7_n31, aluBoi_aluBoi_shft_SLL_sll_7_n30,
         aluBoi_aluBoi_shft_SLL_sll_7_n29, aluBoi_aluBoi_shft_SLL_sll_7_n28,
         aluBoi_aluBoi_shft_SLL_sll_7_n27, aluBoi_aluBoi_shft_SLL_sll_7_n26,
         aluBoi_aluBoi_shft_SLL_sll_7_n25, aluBoi_aluBoi_shft_SLL_sll_7_n24,
         aluBoi_aluBoi_shft_SLL_sll_7_n23, aluBoi_aluBoi_shft_SLL_sll_7_n22,
         aluBoi_aluBoi_shft_SLL_sll_7_n21, aluBoi_aluBoi_shft_SLL_sll_7_n20,
         aluBoi_aluBoi_shft_SLL_sll_7_n19, aluBoi_aluBoi_shft_SLL_sll_7_n18,
         aluBoi_aluBoi_shft_SLL_sll_7_n17, aluBoi_aluBoi_shft_SLL_sll_7_n16,
         aluBoi_aluBoi_shft_SLL_sll_7_n15, aluBoi_aluBoi_shft_SLL_sll_7_n14,
         aluBoi_aluBoi_shft_SLL_sll_7_n13, aluBoi_aluBoi_shft_SLL_sll_7_n12,
         aluBoi_aluBoi_shft_SLL_sll_7_n11, aluBoi_aluBoi_shft_SLL_sll_7_n10,
         aluBoi_aluBoi_shft_SLL_sll_7_n9, aluBoi_aluBoi_shft_SLL_sll_7_n8,
         aluBoi_aluBoi_shft_SLL_sll_7_n7, aluBoi_aluBoi_shft_SLL_sll_7_n6,
         aluBoi_aluBoi_shft_SLL_sll_7_n5, aluBoi_aluBoi_shft_SLL_sll_7_n4,
         aluBoi_aluBoi_shft_SLL_sll_7_n3, aluBoi_aluBoi_shft_SLL_sll_7_n2,
         aluBoi_aluBoi_shft_SLL_sll_7_n1,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__8_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__9_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__10_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__11_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__12_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__13_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__14_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__15_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__16_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__17_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__18_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__19_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__20_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__21_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__22_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__23_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__24_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__25_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__26_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__27_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__28_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__29_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__30_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__31_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__0_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__1_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__2_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__3_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__4_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__5_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__6_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__7_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__8_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__9_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__10_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__11_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__12_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__13_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__14_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__15_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__16_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__17_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__18_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__19_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__20_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__21_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__22_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__23_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__24_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__25_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__26_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__27_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__28_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__29_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__30_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__31_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__0_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__1_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__2_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__3_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__4_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__5_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__6_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__7_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__8_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__9_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__10_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__11_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__12_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__13_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__14_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__15_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__16_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__17_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__18_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__19_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__20_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__21_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__22_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__23_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__24_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__25_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__26_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__27_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__28_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__29_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__30_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__31_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__0_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__1_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__2_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__3_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__4_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__5_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__6_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__7_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__8_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__9_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__10_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__11_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__12_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__13_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__14_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__15_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__16_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__17_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__18_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__19_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__20_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__21_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__22_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__23_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__24_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__25_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__26_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__27_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__28_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__29_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__30_,
         aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__31_;
  wire   [4:0] aluRw;
  wire   [15:7] aluPC8;
  wire   [2:0] aluBoi_multOut;
  wire   [31:0] aluBoi_aluBoi_shft_sraout;
  wire   [31:0] aluBoi_aluBoi_shft_srlout;
  wire   [31:0] aluBoi_aluBoi_shft_sllout;
  wire   [59:0] aluBoi_multBoi_temppp;
  assign daluKill = difHold;
  assign didHold = difHold;

  DFFR_X1 aluBoi_aluReg_75__regBoi_curData_reg ( .D(n4876), .CK(clk), .RN(
        n6884), .Q(daddr[31]), .QN(n5328) );
  DFFR_X1 idBoi_reggal_30__regBoi_curData_reg ( .D(n4874), .CK(clk), .RN(n6921), .Q(didMult) );
  DFFR_X1 ifBoi_reglol_63__regBoi_curData_reg ( .D(n13607), .CK(clk), .RN(
        n6898), .Q(ifInst[31]) );
  DFFR_X1 ifBoi_reglol_61__regBoi_curData_reg ( .D(n13605), .CK(clk), .RN(
        n6898), .Q(ifInst[29]) );
  DFFR_X1 ifBoi_reglol_58__regBoi_curData_reg ( .D(n13602), .CK(clk), .RN(
        n6898), .Q(ifInst[26]) );
  DFFR_X1 ifBoi_reglol_57__regBoi_curData_reg ( .D(n13601), .CK(clk), .RN(
        n6876), .Q(n5313), .QN(n5354) );
  DFFR_X1 ifBoi_reglol_56__regBoi_curData_reg ( .D(n13600), .CK(clk), .RN(
        n6898), .Q(ifInst[24]) );
  DFFR_X1 ifBoi_reglol_55__regBoi_curData_reg ( .D(n13599), .CK(clk), .RN(
        n6876), .Q(ifInst[23]) );
  DFFR_X1 ifBoi_reglol_54__regBoi_curData_reg ( .D(n13598), .CK(clk), .RN(
        n6898), .Q(ifInst[22]) );
  DFFR_X1 ifBoi_reglol_53__regBoi_curData_reg ( .D(n13597), .CK(clk), .RN(
        n6876), .Q(ifInst[21]) );
  DFFR_X1 idBoi_reggal_9__regBoi_curData_reg ( .D(n4841), .CK(clk), .RN(n6896), 
        .Q(aluBoi_imm32w_9_) );
  DFFR_X1 idBoi_reggal_7__regBoi_curData_reg ( .D(n4837), .CK(clk), .RN(n6895), 
        .Q(aluBoi_imm32w_7_) );
  DFFR_X1 idBoi_reggal_74__regBoi_curData_reg ( .D(n4834), .CK(clk), .RN(n6894), .Q(idOut_74_), .QN(n5594) );
  DFFR_X1 idBoi_reggal_72__regBoi_curData_reg ( .D(n4833), .CK(clk), .RN(n6894), .Q(idOut_72_), .QN(n5592) );
  DFFR_X1 idBoi_reggal_5__regBoi_curData_reg ( .D(n4832), .CK(clk), .RN(n6894), 
        .Q(aluBoi_imm32w_5_) );
  DFFR_X1 idBoi_reggal_38__regBoi_curData_reg ( .D(n4830), .CK(clk), .RN(n6893), .Q(idOut_38_) );
  DFFR_X1 idBoi_reggal_34__regBoi_curData_reg ( .D(n4829), .CK(clk), .RN(n6893), .Q(idOut_34_) );
  DFFR_X1 idBoi_reggal_32__regBoi_curData_reg ( .D(n4828), .CK(clk), .RN(n6849), .Q(idOut_32_), .QN(n5522) );
  DFFR_X1 idBoi_reggal_27__regBoi_curData_reg ( .D(n4827), .CK(clk), .RN(n6848), .Q(aluifJRflag), .QN(n5476) );
  DFFR_X1 idBoi_reggal_25__regBoi_curData_reg ( .D(n4826), .CK(clk), .RN(n6845), .Q(idOut_25_), .QN(n5472) );
  DFFR_X1 idBoi_reggal_17__regBoi_curData_reg ( .D(n4825), .CK(clk), .RN(n6882), .Q(idOut_17_), .QN(n5620) );
  DFFR_X1 idBoi_reggal_15__regBoi_curData_reg ( .D(n4824), .CK(clk), .RN(n6882), .Q(aluBoi_imm32w_15_) );
  DFFR_X1 idBoi_reggal_13__regBoi_curData_reg ( .D(n4823), .CK(clk), .RN(n6882), .Q(aluBoi_imm32w_13_) );
  DFFR_X1 idBoi_reggal_11__regBoi_curData_reg ( .D(n4822), .CK(clk), .RN(n6882), .Q(aluBoi_imm32w_11_) );
  DFFR_X1 idBoi_reggal_10__regBoi_curData_reg ( .D(n4820), .CK(clk), .RN(n6892), .Q(aluBoi_imm32w_10_) );
  DFFR_X1 idBoi_reggal_12__regBoi_curData_reg ( .D(n4819), .CK(clk), .RN(n6865), .Q(aluBoi_imm32w_12_) );
  DFFR_X1 idBoi_reggal_14__regBoi_curData_reg ( .D(n4818), .CK(clk), .RN(n6861), .Q(aluBoi_imm32w_14_) );
  DFFR_X1 idBoi_reggal_26__regBoi_curData_reg ( .D(n4816), .CK(clk), .RN(n6881), .Q(idOut_26_) );
  DFFR_X1 idBoi_reggal_31__regBoi_curData_reg ( .D(n4814), .CK(clk), .RN(n6881), .Q(idOut_31_), .QN(n5676) );
  DFFR_X1 idBoi_reggal_33__regBoi_curData_reg ( .D(n4813), .CK(clk), .RN(n6881), .Q(idOut_33_), .QN(n5556) );
  DFFR_X1 idBoi_reggal_6__regBoi_curData_reg ( .D(n13612), .CK(clk), .RN(n6879), .Q(aluBoi_imm32w_6_) );
  DFFR_X1 idBoi_reggal_71__regBoi_curData_reg ( .D(n4810), .CK(clk), .RN(n6879), .Q(idOut_71_), .QN(n5591) );
  DFFR_X1 idBoi_reggal_73__regBoi_curData_reg ( .D(n4809), .CK(clk), .RN(n6879), .Q(idOut_73_), .QN(n5593) );
  DFFR_X1 idBoi_reggal_75__regBoi_curData_reg ( .D(n4808), .CK(clk), .RN(n6879), .Q(idOut_75_), .QN(n5595) );
  DFFR_X1 idBoi_reggal_8__regBoi_curData_reg ( .D(n4802), .CK(clk), .RN(n6878), 
        .Q(aluBoi_imm32w_8_) );
  DFFR_X1 aluBoi_aluReg_38__regBoi_curData_reg ( .D(n13657), .CK(clk), .RN(
        n6889), .Q(dwData[31]) );
  DFFR_X1 aluBoi_aluReg_4__regBoi_curData_reg ( .D(n4794), .CK(clk), .RN(n6885), .Q(dSize[1]), .QN(n5353) );
  DFFR_X1 aluBoi_aluReg_6__regBoi_curData_reg ( .D(n13663), .CK(clk), .RN(
        n6884), .Q(dWr) );
  DFFR_X1 idBoi_reggal_23__regBoi_curData_reg ( .D(n13608), .CK(clk), .RN(
        n6852), .Q(idOut_23_) );
  DFFR_X1 idBoi_reggal_20__regBoi_curData_reg ( .D(n4790), .CK(clk), .RN(n6881), .Q(idOut_20_), .QN(n5716) );
  DFFR_X1 idBoi_reggal_19__regBoi_curData_reg ( .D(n4789), .CK(clk), .RN(n6881), .Q(idOut_19_), .QN(n5715) );
  DFFR_X1 idBoi_reggal_18__regBoi_curData_reg ( .D(n4788), .CK(clk), .RN(n6929), .Q(idOut_18_), .QN(n5391) );
  DFFR_X1 idBoi_reggal_35__regBoi_curData_reg ( .D(n4786), .CK(clk), .RN(n6881), .Q(idRegWr) );
  DFFR_X1 aluBoi_aluReg_0__regBoi_curData_reg ( .D(n13662), .CK(clk), .RN(
        n6887), .Q(aluRegWrOut) );
  DFFR_X1 idBoi_reggal_22__regBoi_curData_reg ( .D(n4784), .CK(clk), .RN(n6881), .Q(idOut_22_), .QN(n5345) );
  DFFR_X1 idBoi_reggal_24__regBoi_curData_reg ( .D(n4783), .CK(clk), .RN(n6881), .Q(idOut_24_) );
  DFFR_X1 idBoi_reggal_21__regBoi_curData_reg ( .D(n4782), .CK(clk), .RN(n6940), .Q(idOut_21_), .QN(n5363) );
  DFFR_X1 aluBoi_aluReg_7__regBoi_curData_reg ( .D(n13658), .CK(clk), .RN(
        n6891), .Q(dwData[0]) );
  DFFR_X1 aluBoi_aluReg_8__regBoi_curData_reg ( .D(n13659), .CK(clk), .RN(
        n6883), .Q(dwData[1]) );
  DFFR_X1 aluBoi_aluReg_46__regBoi_curData_reg ( .D(n4777), .CK(clk), .RN(
        n6885), .Q(daddr[2]) );
  DFFR_X1 aluBoi_aluReg_9__regBoi_curData_reg ( .D(n13660), .CK(clk), .RN(
        n6892), .Q(dwData[2]) );
  DFFR_X1 aluBoi_aluReg_47__regBoi_curData_reg ( .D(n4775), .CK(clk), .RN(
        n6889), .Q(daddr[3]) );
  DFFR_X1 aluBoi_aluReg_10__regBoi_curData_reg ( .D(n13629), .CK(clk), .RN(
        n6888), .Q(dwData[3]) );
  DFFR_X1 aluBoi_aluReg_36__regBoi_curData_reg ( .D(n13655), .CK(clk), .RN(
        n6889), .Q(dwData[29]) );
  DFFR_X1 aluBoi_aluReg_74__regBoi_curData_reg ( .D(n4771), .CK(clk), .RN(
        n6890), .Q(daddr[30]), .QN(n5321) );
  DFFR_X1 aluBoi_aluReg_37__regBoi_curData_reg ( .D(n13656), .CK(clk), .RN(
        n6886), .Q(dwData[30]) );
  DFFR_X1 aluBoi_aluReg_33__regBoi_curData_reg ( .D(n13652), .CK(clk), .RN(
        n6886), .Q(dwData[26]) );
  DFFR_X1 aluBoi_aluReg_34__regBoi_curData_reg ( .D(n13653), .CK(clk), .RN(
        n6889), .Q(dwData[27]) );
  DFFR_X1 aluBoi_aluReg_72__regBoi_curData_reg ( .D(n4765), .CK(clk), .RN(
        n6890), .Q(daddr[28]), .QN(n5320) );
  DFFR_X1 aluBoi_aluReg_35__regBoi_curData_reg ( .D(n13654), .CK(clk), .RN(
        n6886), .Q(dwData[28]) );
  DFFR_X1 aluBoi_aluReg_68__regBoi_curData_reg ( .D(n4763), .CK(clk), .RN(
        n6884), .Q(daddr[24]), .QN(n5325) );
  DFFR_X1 aluBoi_aluReg_31__regBoi_curData_reg ( .D(n13650), .CK(clk), .RN(
        n6886), .Q(dwData[24]) );
  DFFR_X1 aluBoi_aluReg_69__regBoi_curData_reg ( .D(n4761), .CK(clk), .RN(
        n6890), .Q(daddr[25]), .QN(n5326) );
  DFFR_X1 aluBoi_aluReg_32__regBoi_curData_reg ( .D(n13651), .CK(clk), .RN(
        n6889), .Q(dwData[25]) );
  DFFR_X1 aluBoi_aluReg_67__regBoi_curData_reg ( .D(n4759), .CK(clk), .RN(
        n6890), .Q(daddr[23]), .QN(n5324) );
  DFFR_X1 aluBoi_aluReg_30__regBoi_curData_reg ( .D(n13649), .CK(clk), .RN(
        n6888), .Q(dwData[23]) );
  DFFR_X1 aluBoi_aluReg_66__regBoi_curData_reg ( .D(n4757), .CK(clk), .RN(
        n6884), .Q(daddr[22]), .QN(n5503) );
  DFFR_X1 aluBoi_aluReg_29__regBoi_curData_reg ( .D(n13648), .CK(clk), .RN(
        n6888), .Q(dwData[22]) );
  DFFR_X1 aluBoi_aluReg_65__regBoi_curData_reg ( .D(n4755), .CK(clk), .RN(
        n6890), .Q(daddr[21]), .QN(n5502) );
  DFFR_X1 aluBoi_aluReg_28__regBoi_curData_reg ( .D(n13647), .CK(clk), .RN(
        n6886), .Q(dwData[21]) );
  DFFR_X1 aluBoi_aluReg_64__regBoi_curData_reg ( .D(n4753), .CK(clk), .RN(
        n6884), .Q(daddr[20]), .QN(n5501) );
  DFFR_X1 aluBoi_aluReg_23__regBoi_curData_reg ( .D(n13642), .CK(clk), .RN(
        n6888), .Q(dwData[16]) );
  DFFR_X1 aluBoi_aluReg_61__regBoi_curData_reg ( .D(n4750), .CK(clk), .RN(
        n6890), .Q(daddr[17]), .QN(n5499) );
  DFFR_X1 aluBoi_aluReg_24__regBoi_curData_reg ( .D(n13643), .CK(clk), .RN(
        n6886), .Q(dwData[17]) );
  DFFR_X1 aluBoi_aluReg_62__regBoi_curData_reg ( .D(n4748), .CK(clk), .RN(
        n6884), .Q(daddr[18]), .QN(n5500) );
  DFFR_X1 aluBoi_aluReg_25__regBoi_curData_reg ( .D(n13644), .CK(clk), .RN(
        n6888), .Q(dwData[18]) );
  DFFR_X1 aluBoi_aluReg_18__regBoi_curData_reg ( .D(n13637), .CK(clk), .RN(
        n6888), .Q(dwData[11]) );
  DFFR_X1 aluBoi_aluReg_19__regBoi_curData_reg ( .D(n13638), .CK(clk), .RN(
        n6886), .Q(dwData[12]) );
  DFFR_X1 aluBoi_aluReg_20__regBoi_curData_reg ( .D(n13639), .CK(clk), .RN(
        n6886), .Q(dwData[13]) );
  DFFR_X1 aluBoi_aluReg_50__regBoi_curData_reg ( .D(n4738), .CK(clk), .RN(
        n6889), .Q(daddr[6]) );
  DFFR_X1 aluBoi_aluReg_13__regBoi_curData_reg ( .D(n13632), .CK(clk), .RN(
        n6887), .Q(dwData[6]) );
  DFFR_X1 aluBoi_aluReg_51__regBoi_curData_reg ( .D(n4736), .CK(clk), .RN(
        n6885), .Q(daddr[7]) );
  DFFR_X1 aluBoi_aluReg_14__regBoi_curData_reg ( .D(n13633), .CK(clk), .RN(
        n6888), .Q(dwData[7]) );
  DFFR_X1 aluBoi_aluReg_48__regBoi_curData_reg ( .D(n4733), .CK(clk), .RN(
        n6885), .Q(daddr[4]) );
  DFFR_X1 aluBoi_aluReg_11__regBoi_curData_reg ( .D(n13630), .CK(clk), .RN(
        n6887), .Q(dwData[4]) );
  DFFR_X1 aluBoi_aluReg_15__regBoi_curData_reg ( .D(n13634), .CK(clk), .RN(
        n6887), .Q(dwData[8]) );
  DFFR_X1 aluBoi_aluReg_49__regBoi_curData_reg ( .D(n4729), .CK(clk), .RN(
        n6889), .Q(daddr[5]) );
  DFFR_X1 aluBoi_aluReg_12__regBoi_curData_reg ( .D(n13631), .CK(clk), .RN(
        n6888), .Q(dwData[5]) );
  DFFR_X1 aluBoi_aluReg_16__regBoi_curData_reg ( .D(n13635), .CK(clk), .RN(
        n6888), .Q(dwData[9]) );
  DFFR_X1 aluBoi_aluReg_17__regBoi_curData_reg ( .D(n13636), .CK(clk), .RN(
        n6886), .Q(dwData[10]) );
  DFFR_X1 aluBoi_aluReg_21__regBoi_curData_reg ( .D(n13640), .CK(clk), .RN(
        n6888), .Q(dwData[14]) );
  DFFR_X1 aluBoi_aluReg_22__regBoi_curData_reg ( .D(n13641), .CK(clk), .RN(
        n6886), .Q(dwData[15]) );
  DFFR_X1 aluBoi_aluReg_26__regBoi_curData_reg ( .D(n13645), .CK(clk), .RN(
        n6886), .Q(dwData[19]) );
  DFFR_X1 aluBoi_aluReg_27__regBoi_curData_reg ( .D(n13646), .CK(clk), .RN(
        n6888), .Q(dwData[20]) );
  DFFR_X1 idBoi_reggal_28__regBoi_curData_reg ( .D(n4719), .CK(clk), .RN(n6881), .Q(idOut_28_), .QN(n5621) );
  DFFR_X1 aluBoi_aluReg_5__regBoi_curData_reg ( .D(n4718), .CK(clk), .RN(n6890), .Q(aluDExtOp), .QN(n5384) );
  DFFR_X1 idBoi_reggal_16__regBoi_curData_reg ( .D(n4717), .CK(clk), .RN(n6842), .Q(idOut_16_), .QN(n5619) );
  DFFR_X1 aluBoi_aluReg_3__regBoi_curData_reg ( .D(n4716), .CK(clk), .RN(n6889), .Q(dSize[0]), .QN(n5318) );
  DFFR_X1 idBoi_reggal_36__regBoi_curData_reg ( .D(n4715), .CK(clk), .RN(n6893), .QN(n5583) );
  DFFR_X1 aluBoi_aluReg_1__regBoi_curData_reg ( .D(n4714), .CK(clk), .RN(n6888), .Q(aluMem2Reg), .QN(n5519) );
  DFFR_X1 ifBoi_reglol_64__regBoi_curData_reg ( .D(n4712), .CK(clk), .RN(n6884), .Q(ifOut_64_) );
  DFFR_X1 idBoi_reggal_86__regBoi_curData_reg ( .D(n4711), .CK(clk), .RN(n6878), .Q(idOut_86_) );
  DFFR_X1 ifBoi_reglol_0__regBoi_curData_reg ( .D(n4710), .CK(clk), .RN(n6878), 
        .Q(ifOut_0_) );
  DFFR_X1 idBoi_reggal_39__regBoi_curData_reg ( .D(n4709), .CK(clk), .RN(n6881), .Q(idOut_39_), .QN(n5622) );
  DFFR_X1 idBoi_reggal_87__regBoi_curData_reg ( .D(n4706), .CK(clk), .RN(n6895), .Q(idOut_87_) );
  DFFR_X1 ifBoi_reglol_1__regBoi_curData_reg ( .D(n4705), .CK(clk), .RN(n6896), 
        .Q(ifOut_1_) );
  DFFR_X1 idBoi_reggal_40__regBoi_curData_reg ( .D(n4704), .CK(clk), .RN(n6880), .Q(idOut_40_), .QN(n5623) );
  DFFR_X1 ifBoi_reglol_2__regBoi_curData_reg ( .D(n4700), .CK(clk), .RN(n6877), 
        .Q(ifOut_2_), .QN(n5610) );
  DFFR_X1 idBoi_reggal_41__regBoi_curData_reg ( .D(n4699), .CK(clk), .RN(n6893), .Q(idOut_41_), .QN(n5624) );
  DFFR_X1 ifBoi_reglol_3__regBoi_curData_reg ( .D(n4697), .CK(clk), .RN(n6897), 
        .Q(ifOut_3_) );
  DFFR_X1 idBoi_reggal_42__regBoi_curData_reg ( .D(n4696), .CK(clk), .RN(n6880), .Q(idOut_42_), .QN(n5625) );
  DFFR_X1 ifBoi_reglol_67__regBoi_curData_reg ( .D(n4695), .CK(clk), .RN(n6898), .Q(ifOut_67_) );
  DFFR_X1 idBoi_reggal_89__regBoi_curData_reg ( .D(n13623), .CK(clk), .RN(
        n6895), .Q(idOut_89_) );
  DFFR_X1 ifBoi_reglol_4__regBoi_curData_reg ( .D(n4692), .CK(clk), .RN(n6876), 
        .Q(ifOut_4_) );
  DFFR_X1 idBoi_reggal_43__regBoi_curData_reg ( .D(n4691), .CK(clk), .RN(n6893), .Q(idOut_43_), .QN(n5626) );
  DFFR_X1 idBoi_reggal_90__regBoi_curData_reg ( .D(n4689), .CK(clk), .RN(n6895), .Q(idOut_90_) );
  DFFR_X1 ifBoi_reglol_5__regBoi_curData_reg ( .D(n4687), .CK(clk), .RN(n6898), 
        .Q(ifOut_5_) );
  DFFR_X1 idBoi_reggal_44__regBoi_curData_reg ( .D(n4686), .CK(clk), .RN(n6880), .Q(idOut_44_), .QN(n5627) );
  DFFR_X1 ifBoi_reglol_69__regBoi_curData_reg ( .D(n4685), .CK(clk), .RN(n6898), .Q(ifOut_69_) );
  DFFR_X1 idBoi_reggal_91__regBoi_curData_reg ( .D(n13624), .CK(clk), .RN(
        n6878), .Q(idOut_91_) );
  DFFR_X1 ifBoi_reglol_6__regBoi_curData_reg ( .D(n4682), .CK(clk), .RN(n6941), 
        .Q(ifOut_6_), .QN(n5609) );
  DFFR_X1 idBoi_reggal_45__regBoi_curData_reg ( .D(n4681), .CK(clk), .RN(n6893), .Q(idOut_45_), .QN(n5628) );
  DFFR_X1 idBoi_reggal_92__regBoi_curData_reg ( .D(n4679), .CK(clk), .RN(n6895), .Q(idOut_92_) );
  DFFR_X1 ifBoi_reglol_7__regBoi_curData_reg ( .D(n4677), .CK(clk), .RN(n6899), 
        .Q(ifOut_7_) );
  DFFR_X1 idBoi_reggal_46__regBoi_curData_reg ( .D(n4676), .CK(clk), .RN(n6880), .Q(idOut_46_) );
  DFFR_X1 ifBoi_reglol_71__regBoi_curData_reg ( .D(n4675), .CK(clk), .RN(n6935), .Q(ifOut_71_) );
  DFFR_X1 idBoi_reggal_93__regBoi_curData_reg ( .D(n13625), .CK(clk), .RN(
        n6878), .Q(idOut_93_) );
  DFFR_X1 ifBoi_reglol_8__regBoi_curData_reg ( .D(n4672), .CK(clk), .RN(n6875), 
        .Q(ifOut_8_), .QN(n5608) );
  DFFR_X1 idBoi_reggal_47__regBoi_curData_reg ( .D(n4671), .CK(clk), .RN(n6893), .Q(idOut_47_) );
  DFFR_X1 idBoi_reggal_94__regBoi_curData_reg ( .D(n4669), .CK(clk), .RN(n6895), .Q(idOut_94_) );
  DFFR_X1 ifBoi_reglol_9__regBoi_curData_reg ( .D(n4667), .CK(clk), .RN(n6900), 
        .Q(ifOut_9_) );
  DFFR_X1 idBoi_reggal_48__regBoi_curData_reg ( .D(n13610), .CK(clk), .RN(
        n6880), .Q(idOut_48_) );
  DFFR_X1 ifBoi_reglol_73__regBoi_curData_reg ( .D(n4665), .CK(clk), .RN(n6927), .Q(ifOut_73_) );
  DFFR_X1 idBoi_reggal_95__regBoi_curData_reg ( .D(n13626), .CK(clk), .RN(
        n6878), .Q(idOut_95_) );
  DFFR_X1 idBoi_reggal_96__regBoi_curData_reg ( .D(n4661), .CK(clk), .RN(n6895), .Q(idOut_96_) );
  DFFR_X1 ifBoi_reglol_10__regBoi_curData_reg ( .D(n4660), .CK(clk), .RN(n6896), .Q(ifOut_10_), .QN(n5607) );
  DFFR_X1 idBoi_reggal_49__regBoi_curData_reg ( .D(n13611), .CK(clk), .RN(
        n6893), .Q(idOut_49_) );
  DFFR_X1 ifBoi_reglol_11__regBoi_curData_reg ( .D(n4657), .CK(clk), .RN(n6878), .Q(ifOut_11_) );
  DFFR_X1 idBoi_reggal_50__regBoi_curData_reg ( .D(n4656), .CK(clk), .RN(n6893), .Q(idOut_50_) );
  DFFR_X1 ifBoi_reglol_75__regBoi_curData_reg ( .D(n4655), .CK(clk), .RN(n6881), .Q(ifOut_75_) );
  DFFR_X1 idBoi_reggal_97__regBoi_curData_reg ( .D(n13627), .CK(clk), .RN(
        n6878), .Q(idOut_97_) );
  DFFR_X1 ifBoi_reglol_76__regBoi_curData_reg ( .D(n4652), .CK(clk), .RN(n6899), .Q(ifOut_76_) );
  DFFR_X1 idBoi_reggal_98__regBoi_curData_reg ( .D(n4651), .CK(clk), .RN(n6895), .Q(idOut_98_) );
  DFFR_X1 ifBoi_reglol_12__regBoi_curData_reg ( .D(n4650), .CK(clk), .RN(n6896), .Q(ifOut_12_) );
  DFFR_X1 idBoi_reggal_51__regBoi_curData_reg ( .D(n4649), .CK(clk), .RN(n6880), .Q(idOut_51_) );
  DFFR_X1 ifBoi_reglol_13__regBoi_curData_reg ( .D(n4647), .CK(clk), .RN(n6878), .Q(ifOut_13_), .QN(n5606) );
  DFFR_X1 idBoi_reggal_52__regBoi_curData_reg ( .D(n4646), .CK(clk), .RN(n6893), .Q(idOut_52_) );
  DFFR_X1 ifBoi_reglol_77__regBoi_curData_reg ( .D(n4645), .CK(clk), .RN(n6859), .Q(ifOut_77_) );
  DFFR_X1 idBoi_reggal_99__regBoi_curData_reg ( .D(n13628), .CK(clk), .RN(
        n6878), .Q(idOut_99_) );
  DFFR_X1 ifBoi_reglol_78__regBoi_curData_reg ( .D(n4642), .CK(clk), .RN(n6899), .Q(ifOut_78_) );
  DFFR_X1 idBoi_reggal_100__regBoi_curData_reg ( .D(n4641), .CK(clk), .RN(
        n6892), .Q(idOut_100_) );
  DFFR_X1 ifBoi_reglol_14__regBoi_curData_reg ( .D(n4640), .CK(clk), .RN(n6896), .Q(ifOut_14_) );
  DFFR_X1 idBoi_reggal_53__regBoi_curData_reg ( .D(n4639), .CK(clk), .RN(n6880), .Q(idOut_53_) );
  DFFR_X1 ifBoi_reglol_15__regBoi_curData_reg ( .D(n4637), .CK(clk), .RN(n6877), .Q(ifOut_15_), .QN(n5605) );
  DFFR_X1 idBoi_reggal_54__regBoi_curData_reg ( .D(n4636), .CK(clk), .RN(n6893), .Q(idOut_54_) );
  DFFR_X1 ifBoi_reglol_79__regBoi_curData_reg ( .D(n4635), .CK(clk), .RN(n6914), .Q(ifOut_79_) );
  DFFR_X1 idBoi_reggal_101__regBoi_curData_reg ( .D(n13609), .CK(clk), .RN(
        n6883), .Q(idOut_101_) );
  DFFR_X1 ifBoi_reglol_80__regBoi_curData_reg ( .D(n4632), .CK(clk), .RN(n6875), .Q(ifOut_80_) );
  DFFR_X1 idBoi_reggal_102__regBoi_curData_reg ( .D(n4631), .CK(clk), .RN(
        n6892), .Q(idOut_102_), .QN(n5512) );
  DFFR_X1 ifBoi_reglol_16__regBoi_curData_reg ( .D(n4630), .CK(clk), .RN(n6896), .Q(ifOut_16_) );
  DFFR_X1 idBoi_reggal_55__regBoi_curData_reg ( .D(n4629), .CK(clk), .RN(n6880), .Q(idOut_55_), .QN(n5629) );
  DFFR_X1 ifBoi_reglol_17__regBoi_curData_reg ( .D(n4627), .CK(clk), .RN(n6877), .Q(ifOut_17_), .QN(n5604) );
  DFFR_X1 idBoi_reggal_56__regBoi_curData_reg ( .D(n4626), .CK(clk), .RN(n6894), .Q(idOut_56_), .QN(n5630) );
  DFFR_X1 ifBoi_reglol_81__regBoi_curData_reg ( .D(n4625), .CK(clk), .RN(n6899), .Q(ifOut_81_) );
  DFFR_X1 idBoi_reggal_103__regBoi_curData_reg ( .D(n4624), .CK(clk), .RN(
        n6882), .Q(idOut_103_), .QN(n5523) );
  DFFR_X1 ifBoi_reglol_82__regBoi_curData_reg ( .D(n4622), .CK(clk), .RN(n6875), .Q(ifOut_82_) );
  DFFR_X1 idBoi_reggal_104__regBoi_curData_reg ( .D(n4621), .CK(clk), .RN(
        n6892), .Q(idOut_104_), .QN(n5486) );
  DFFR_X1 ifBoi_reglol_18__regBoi_curData_reg ( .D(n4620), .CK(clk), .RN(n6896), .Q(ifOut_18_) );
  DFFR_X1 idBoi_reggal_57__regBoi_curData_reg ( .D(n4619), .CK(clk), .RN(n6880), .Q(idOut_57_), .QN(n5631) );
  DFFR_X1 ifBoi_reglol_19__regBoi_curData_reg ( .D(n4617), .CK(clk), .RN(n6877), .Q(ifOut_19_), .QN(n5603) );
  DFFR_X1 idBoi_reggal_58__regBoi_curData_reg ( .D(n4616), .CK(clk), .RN(n6894), .Q(idOut_58_), .QN(n5632) );
  DFFR_X1 ifBoi_reglol_83__regBoi_curData_reg ( .D(n4615), .CK(clk), .RN(n6899), .Q(ifOut_83_) );
  DFFR_X1 idBoi_reggal_105__regBoi_curData_reg ( .D(n4614), .CK(clk), .RN(
        n6882), .Q(idOut_105_), .QN(n5518) );
  DFFR_X1 ifBoi_reglol_84__regBoi_curData_reg ( .D(n4612), .CK(clk), .RN(n6875), .Q(ifOut_84_) );
  DFFR_X1 idBoi_reggal_106__regBoi_curData_reg ( .D(n4611), .CK(clk), .RN(
        n6892), .Q(idOut_106_), .QN(n5513) );
  DFFR_X1 ifBoi_reglol_20__regBoi_curData_reg ( .D(n4610), .CK(clk), .RN(n6877), .Q(ifOut_20_) );
  DFFR_X1 idBoi_reggal_59__regBoi_curData_reg ( .D(n4609), .CK(clk), .RN(n6880), .Q(idOut_59_), .QN(n5633) );
  DFFR_X1 ifBoi_reglol_21__regBoi_curData_reg ( .D(n4607), .CK(clk), .RN(n6896), .Q(ifOut_21_), .QN(n5602) );
  DFFR_X1 idBoi_reggal_60__regBoi_curData_reg ( .D(n4606), .CK(clk), .RN(n6880), .Q(idOut_60_), .QN(n5634) );
  DFFR_X1 ifBoi_reglol_85__regBoi_curData_reg ( .D(n4605), .CK(clk), .RN(n6899), .Q(ifOut_85_) );
  DFFR_X1 idBoi_reggal_107__regBoi_curData_reg ( .D(n4604), .CK(clk), .RN(
        n6882), .Q(idOut_107_), .QN(n5504) );
  DFFR_X1 ifBoi_reglol_86__regBoi_curData_reg ( .D(n4602), .CK(clk), .RN(n6875), .Q(ifOut_86_) );
  DFFR_X1 idBoi_reggal_108__regBoi_curData_reg ( .D(n4601), .CK(clk), .RN(
        n6892), .Q(idOut_108_), .QN(n5514) );
  DFFR_X1 ifBoi_reglol_22__regBoi_curData_reg ( .D(n4600), .CK(clk), .RN(n6877), .Q(ifOut_22_) );
  DFFR_X1 idBoi_reggal_61__regBoi_curData_reg ( .D(n4599), .CK(clk), .RN(n6894), .Q(idOut_61_), .QN(n5635) );
  DFFR_X1 ifBoi_reglol_23__regBoi_curData_reg ( .D(n4597), .CK(clk), .RN(n6896), .Q(ifOut_23_) );
  DFFR_X1 idBoi_reggal_62__regBoi_curData_reg ( .D(n4596), .CK(clk), .RN(n6879), .Q(idOut_62_), .QN(n5636) );
  DFFR_X1 ifBoi_reglol_87__regBoi_curData_reg ( .D(n4595), .CK(clk), .RN(n6899), .Q(ifOut_87_) );
  DFFR_X1 idBoi_reggal_109__regBoi_curData_reg ( .D(n4594), .CK(clk), .RN(
        n6882), .Q(idOut_109_), .QN(n5515) );
  DFFR_X1 ifBoi_reglol_88__regBoi_curData_reg ( .D(n4592), .CK(clk), .RN(n6875), .Q(ifOut_88_) );
  DFFR_X1 idBoi_reggal_110__regBoi_curData_reg ( .D(n4591), .CK(clk), .RN(
        n6882), .Q(idOut_110_), .QN(n5524) );
  DFFR_X1 ifBoi_reglol_24__regBoi_curData_reg ( .D(n4590), .CK(clk), .RN(n6877), .Q(ifOut_24_) );
  DFFR_X1 idBoi_reggal_63__regBoi_curData_reg ( .D(n4589), .CK(clk), .RN(n6894), .Q(idOut_63_), .QN(n5611) );
  DFFR_X1 ifBoi_reglol_25__regBoi_curData_reg ( .D(n4587), .CK(clk), .RN(n6896), .Q(ifOut_25_), .QN(n5601) );
  DFFR_X1 idBoi_reggal_64__regBoi_curData_reg ( .D(n4586), .CK(clk), .RN(n6879), .Q(idOut_64_), .QN(n5612) );
  DFFR_X1 ifBoi_reglol_89__regBoi_curData_reg ( .D(n4585), .CK(clk), .RN(n6899), .Q(ifOut_89_) );
  DFFR_X1 idBoi_reggal_111__regBoi_curData_reg ( .D(n4584), .CK(clk), .RN(
        n6892), .Q(idOut_111_), .QN(n5516) );
  DFFR_X1 ifBoi_reglol_90__regBoi_curData_reg ( .D(n4582), .CK(clk), .RN(n6899), .Q(ifOut_90_) );
  DFFR_X1 idBoi_reggal_112__regBoi_curData_reg ( .D(n4581), .CK(clk), .RN(
        n6882), .Q(idOut_112_), .QN(n5505) );
  DFFR_X1 ifBoi_reglol_26__regBoi_curData_reg ( .D(n4580), .CK(clk), .RN(n6877), .Q(ifOut_26_) );
  DFFR_X1 idBoi_reggal_65__regBoi_curData_reg ( .D(n4579), .CK(clk), .RN(n6894), .Q(idOut_65_), .QN(n5613) );
  DFFR_X1 ifBoi_reglol_27__regBoi_curData_reg ( .D(n4577), .CK(clk), .RN(n6896), .Q(ifOut_27_), .QN(n5600) );
  DFFR_X1 idBoi_reggal_66__regBoi_curData_reg ( .D(n4576), .CK(clk), .RN(n6879), .Q(idOut_66_), .QN(n5614) );
  DFFR_X1 ifBoi_reglol_91__regBoi_curData_reg ( .D(n4575), .CK(clk), .RN(n6875), .Q(ifOut_91_) );
  DFFR_X1 idBoi_reggal_113__regBoi_curData_reg ( .D(n4574), .CK(clk), .RN(
        n6892), .Q(idOut_113_), .QN(n5517) );
  DFFR_X1 idBoi_reggal_114__regBoi_curData_reg ( .D(n4571), .CK(clk), .RN(
        n6882), .Q(idOut_114_), .QN(n5462) );
  DFFR_X1 ifBoi_reglol_28__regBoi_curData_reg ( .D(n4570), .CK(clk), .RN(n6877), .Q(ifOut_28_) );
  DFFR_X1 idBoi_reggal_67__regBoi_curData_reg ( .D(n4569), .CK(clk), .RN(n6894), .Q(idOut_67_), .QN(n5615) );
  DFFR_X1 ifBoi_reglol_29__regBoi_curData_reg ( .D(n4567), .CK(clk), .RN(n6896), .Q(ifOut_29_), .QN(n5599) );
  DFFR_X1 idBoi_reggal_68__regBoi_curData_reg ( .D(n4566), .CK(clk), .RN(n6879), .Q(idOut_68_), .QN(n5616) );
  DFFR_X1 ifBoi_reglol_93__regBoi_curData_reg ( .D(n4565), .CK(clk), .RN(n6875), .Q(ifOut_93_), .QN(n5458) );
  DFFR_X1 idBoi_reggal_115__regBoi_curData_reg ( .D(n4564), .CK(clk), .RN(
        n6892), .Q(idOut_115_), .QN(n5350) );
  DFFR_X1 ifBoi_reglol_30__regBoi_curData_reg ( .D(n4562), .CK(clk), .RN(n6897), .Q(ifOut_30_) );
  DFFR_X1 idBoi_reggal_69__regBoi_curData_reg ( .D(n4561), .CK(clk), .RN(n6894), .Q(idOut_69_), .QN(n5617) );
  DFFR_X1 ifBoi_reglol_94__regBoi_curData_reg ( .D(n4560), .CK(clk), .RN(n6899), .Q(ifOut_94_), .QN(n5461) );
  DFFR_X1 idBoi_reggal_116__regBoi_curData_reg ( .D(n4559), .CK(clk), .RN(
        n6882), .Q(idOut_116_), .QN(n5349) );
  DFFR_X1 ifBoi_reglol_31__regBoi_curData_reg ( .D(n4557), .CK(clk), .RN(n6877), .Q(ifOut_31_) );
  DFFR_X1 idBoi_reggal_70__regBoi_curData_reg ( .D(n4556), .CK(clk), .RN(n6894), .Q(idOut_70_), .QN(n5618) );
  DFFR_X1 ifBoi_reglol_95__regBoi_curData_reg ( .D(n4555), .CK(clk), .RN(n6875), .Q(ifOut_95_) );
  DFFR_X1 idBoi_reggal_117__regBoi_curData_reg ( .D(n4554), .CK(clk), .RN(
        n6892), .Q(idOut_117_), .QN(n5554) );
  DFFR_X1 aluBoi_aluReg_76__regBoi_curData_reg ( .D(n4553), .CK(clk), .RN(
        n6891), .QN(n5359) );
  DFFR_X1 aluBoi_aluReg_77__regBoi_curData_reg ( .D(n4552), .CK(clk), .RN(
        n6884), .QN(n5360) );
  DFFR_X1 aluBoi_aluReg_78__regBoi_curData_reg ( .D(n4551), .CK(clk), .RN(
        n6891), .QN(n5361) );
  DFFR_X1 aluBoi_aluReg_79__regBoi_curData_reg ( .D(n4550), .CK(clk), .RN(
        n6884), .QN(n5362) );
  DFFR_X1 aluBoi_aluReg_80__regBoi_curData_reg ( .D(n4549), .CK(clk), .RN(
        n6884), .QN(n5356) );
  DFFR_X1 aluBoi_aluReg_81__regBoi_curData_reg ( .D(n4548), .CK(clk), .RN(
        n6891), .QN(n5357) );
  DFFR_X1 aluBoi_aluReg_82__regBoi_curData_reg ( .D(n4547), .CK(clk), .RN(
        n6883), .QN(n5358) );
  DFFR_X1 aluBoi_aluReg_83__regBoi_curData_reg ( .D(n13664), .CK(clk), .RN(
        n6891), .Q(aluPC8[7]) );
  DFFR_X1 aluBoi_aluReg_84__regBoi_curData_reg ( .D(n13665), .CK(clk), .RN(
        n6883), .Q(aluPC8[8]) );
  DFFR_X1 aluBoi_aluReg_85__regBoi_curData_reg ( .D(n13666), .CK(clk), .RN(
        n6891), .Q(aluPC8[9]) );
  DFFR_X1 aluBoi_aluReg_86__regBoi_curData_reg ( .D(n13667), .CK(clk), .RN(
        n6883), .Q(aluPC8[10]) );
  DFFR_X1 aluBoi_aluReg_87__regBoi_curData_reg ( .D(n13668), .CK(clk), .RN(
        n6891), .Q(aluPC8[11]) );
  DFFR_X1 aluBoi_aluReg_88__regBoi_curData_reg ( .D(n13669), .CK(clk), .RN(
        n6883), .Q(aluPC8[12]) );
  DFFR_X1 aluBoi_aluReg_89__regBoi_curData_reg ( .D(n13670), .CK(clk), .RN(
        n6891), .Q(aluPC8[13]) );
  DFFR_X1 aluBoi_aluReg_90__regBoi_curData_reg ( .D(n13671), .CK(clk), .RN(
        n6891), .Q(aluPC8[14]) );
  DFFR_X1 aluBoi_aluReg_91__regBoi_curData_reg ( .D(n13672), .CK(clk), .RN(
        n6883), .Q(aluPC8[15]) );
  DFFR_X1 aluBoi_aluReg_92__regBoi_curData_reg ( .D(n4537), .CK(clk), .RN(
        n6891), .QN(n5364) );
  DFFR_X1 aluBoi_aluReg_93__regBoi_curData_reg ( .D(n4536), .CK(clk), .RN(
        n6883), .QN(n5365) );
  DFFR_X1 aluBoi_aluReg_94__regBoi_curData_reg ( .D(n4535), .CK(clk), .RN(
        n6891), .QN(n5366) );
  DFFR_X1 aluBoi_aluReg_95__regBoi_curData_reg ( .D(n4534), .CK(clk), .RN(
        n6883), .QN(n5367) );
  DFFR_X1 aluBoi_aluReg_96__regBoi_curData_reg ( .D(n4533), .CK(clk), .RN(
        n6891), .QN(n5368) );
  DFFR_X1 aluBoi_aluReg_97__regBoi_curData_reg ( .D(n4532), .CK(clk), .RN(
        n6883), .QN(n5369) );
  DFFR_X1 aluBoi_aluReg_98__regBoi_curData_reg ( .D(n4531), .CK(clk), .RN(
        n6892), .QN(n5370) );
  DFFR_X1 aluBoi_aluReg_99__regBoi_curData_reg ( .D(n4530), .CK(clk), .RN(
        n6883), .QN(n5371) );
  DFFR_X1 aluBoi_aluReg_100__regBoi_curData_reg ( .D(n4529), .CK(clk), .RN(
        n6887), .QN(n5372) );
  DFFR_X1 aluBoi_aluReg_101__regBoi_curData_reg ( .D(n4528), .CK(clk), .RN(
        n6887), .QN(n5373) );
  DFFR_X1 aluBoi_aluReg_102__regBoi_curData_reg ( .D(n4527), .CK(clk), .RN(
        n6887), .QN(n5329) );
  DFFR_X1 aluBoi_aluReg_103__regBoi_curData_reg ( .D(n4526), .CK(clk), .RN(
        n6887), .QN(n5330) );
  DFFR_X1 aluBoi_aluReg_104__regBoi_curData_reg ( .D(n4525), .CK(clk), .RN(
        n6887), .QN(n5374) );
  DFFR_X1 aluBoi_aluReg_105__regBoi_curData_reg ( .D(n4524), .CK(clk), .RN(
        n6887), .QN(n5375) );
  DFFR_X1 aluBoi_aluReg_106__regBoi_curData_reg ( .D(n4523), .CK(clk), .RN(
        n6887), .QN(n5376) );
  DFFR_X1 aluBoi_aluReg_107__regBoi_curData_reg ( .D(n4522), .CK(clk), .RN(
        n6887), .QN(n5377) );
  DFFR_X1 memBoi_memReg_0__regBoi_curData_reg ( .D(n5898), .CK(clk), .RN(n6875), .Q(wbRwh[0]), .QN(n5511) );
  DFFR_X1 memBoi_memReg_1__regBoi_curData_reg ( .D(aluRw[1]), .CK(clk), .RN(
        n6900), .Q(wbRwh[1]) );
  DFFR_X1 memBoi_memReg_2__regBoi_curData_reg ( .D(aluRw[2]), .CK(clk), .RN(
        n6874), .Q(wbRwh[2]), .QN(n5482) );
  DFFR_X1 memBoi_memReg_3__regBoi_curData_reg ( .D(aluRw[3]), .CK(clk), .RN(
        n6901), .Q(wbRwh[3]) );
  DFFR_X1 memBoi_memReg_4__regBoi_curData_reg ( .D(aluRw[4]), .CK(clk), .RN(
        n6873), .Q(wbRwh[4]) );
  DFFR_X1 memBoi_memReg_5__regBoi_curData_reg ( .D(aluRegWrOut), .CK(clk), 
        .RN(n6901), .Q(wbRegWrh), .QN(n5565) );
  DFFR_X1 memBoi_memReg_6__regBoi_curData_reg ( .D(n4521), .CK(clk), .RN(n6873), .Q(wbBusWh[0]), .QN(n5683) );
  DFFR_X1 regBoiz_regfile_reg_31__31_ ( .D(n4520), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__31_) );
  DFFR_X1 regBoiz_regfile_reg_30__31_ ( .D(n4519), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_30__31_) );
  DFFR_X1 regBoiz_regfile_reg_29__31_ ( .D(n4518), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__31_) );
  DFFR_X1 regBoiz_regfile_reg_28__31_ ( .D(n4517), .CK(clk), .RN(n6879), .Q(
        regBoiz_regfile_28__31_) );
  DFFR_X1 regBoiz_regfile_reg_27__31_ ( .D(n4516), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__31_) );
  DFFR_X1 regBoiz_regfile_reg_26__31_ ( .D(n4515), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__31_) );
  DFFR_X1 regBoiz_regfile_reg_25__31_ ( .D(n4514), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_25__31_) );
  DFFR_X1 regBoiz_regfile_reg_24__31_ ( .D(n4513), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__31_) );
  DFFR_X1 regBoiz_regfile_reg_23__31_ ( .D(n4512), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__31_) );
  DFFR_X1 regBoiz_regfile_reg_22__31_ ( .D(n4511), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_22__31_) );
  DFFR_X1 regBoiz_regfile_reg_21__31_ ( .D(n4510), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__31_) );
  DFFR_X1 regBoiz_regfile_reg_20__31_ ( .D(n4509), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__31_) );
  DFFR_X1 regBoiz_regfile_reg_19__31_ ( .D(n4508), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__31_) );
  DFFR_X1 regBoiz_regfile_reg_18__31_ ( .D(n4507), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__31_) );
  DFFR_X1 regBoiz_regfile_reg_17__31_ ( .D(n4506), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_17__31_) );
  DFFR_X1 regBoiz_regfile_reg_16__31_ ( .D(n4505), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__31_) );
  DFFR_X1 regBoiz_regfile_reg_15__31_ ( .D(n4504), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__31_), .QN(n5598) );
  DFFR_X1 regBoiz_regfile_reg_14__31_ ( .D(n4503), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_14__31_) );
  DFFR_X1 regBoiz_regfile_reg_13__31_ ( .D(n4502), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__31_), .QN(n5597) );
  DFFR_X1 regBoiz_regfile_reg_12__31_ ( .D(n4501), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__31_) );
  DFFR_X1 regBoiz_regfile_reg_11__31_ ( .D(n4500), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_11__31_), .QN(n5570) );
  DFFR_X1 regBoiz_regfile_reg_9__31_ ( .D(n4498), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_9__31_), .QN(n5590) );
  DFFR_X1 regBoiz_regfile_reg_7__31_ ( .D(n4496), .CK(clk), .RN(n6893), .Q(
        regBoiz_regfile_7__31_) );
  DFFR_X1 regBoiz_regfile_reg_6__31_ ( .D(n4495), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__31_) );
  DFFR_X1 regBoiz_regfile_reg_5__31_ ( .D(n4494), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__31_) );
  DFFR_X1 regBoiz_regfile_reg_4__31_ ( .D(n4493), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_4__31_) );
  DFFR_X1 regBoiz_regfile_reg_3__31_ ( .D(n4492), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__31_), .QN(n5576) );
  DFFR_X1 regBoiz_regfile_reg_1__31_ ( .D(n4490), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_1__31_), .QN(n5577) );
  DFFR_X1 regBoiz_regfile_reg_0__31_ ( .D(n4489), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__31_) );
  DFFR_X1 memBoi_memReg_7__regBoi_curData_reg ( .D(n4488), .CK(clk), .RN(n6901), .Q(wbBusWh[1]), .QN(n5670) );
  DFFR_X1 regBoiz_regfile_reg_31__30_ ( .D(n4487), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__30_) );
  DFFR_X1 regBoiz_regfile_reg_30__30_ ( .D(n4486), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__30_) );
  DFFR_X1 regBoiz_regfile_reg_29__30_ ( .D(n4485), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__30_) );
  DFFR_X1 regBoiz_regfile_reg_28__30_ ( .D(n4484), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__30_) );
  DFFR_X1 regBoiz_regfile_reg_27__30_ ( .D(n4483), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__30_) );
  DFFR_X1 regBoiz_regfile_reg_26__30_ ( .D(n4482), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__30_) );
  DFFR_X1 regBoiz_regfile_reg_25__30_ ( .D(n4481), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__30_), .QN(n5759) );
  DFFR_X1 regBoiz_regfile_reg_24__30_ ( .D(n4480), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__30_), .QN(n5760) );
  DFFR_X1 regBoiz_regfile_reg_23__30_ ( .D(n4479), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__30_) );
  DFFR_X1 regBoiz_regfile_reg_22__30_ ( .D(n4478), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__30_) );
  DFFR_X1 regBoiz_regfile_reg_21__30_ ( .D(n4477), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__30_) );
  DFFR_X1 regBoiz_regfile_reg_20__30_ ( .D(n4476), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__30_) );
  DFFR_X1 regBoiz_regfile_reg_19__30_ ( .D(n4475), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__30_) );
  DFFR_X1 regBoiz_regfile_reg_18__30_ ( .D(n4474), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__30_) );
  DFFR_X1 regBoiz_regfile_reg_17__30_ ( .D(n4473), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__30_) );
  DFFR_X1 regBoiz_regfile_reg_16__30_ ( .D(n4472), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__30_) );
  DFFR_X1 regBoiz_regfile_reg_15__30_ ( .D(n4471), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__30_) );
  DFFR_X1 regBoiz_regfile_reg_14__30_ ( .D(n4470), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__30_), .QN(n5408) );
  DFFR_X1 regBoiz_regfile_reg_13__30_ ( .D(n4469), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__30_) );
  DFFR_X1 regBoiz_regfile_reg_12__30_ ( .D(n4468), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__30_), .QN(n5409) );
  DFFR_X1 regBoiz_regfile_reg_11__30_ ( .D(n4467), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__30_) );
  DFFR_X1 regBoiz_regfile_reg_10__30_ ( .D(n4466), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__30_) );
  DFFR_X1 regBoiz_regfile_reg_9__30_ ( .D(n4465), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_9__30_) );
  DFFR_X1 regBoiz_regfile_reg_8__30_ ( .D(n4464), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__30_) );
  DFFR_X1 regBoiz_regfile_reg_7__30_ ( .D(n4463), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__30_) );
  DFFR_X1 regBoiz_regfile_reg_6__30_ ( .D(n4462), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__30_) );
  DFFR_X1 regBoiz_regfile_reg_5__30_ ( .D(n4461), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__30_) );
  DFFR_X1 regBoiz_regfile_reg_4__30_ ( .D(n4460), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__30_) );
  DFFR_X1 regBoiz_regfile_reg_3__30_ ( .D(n4459), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__30_) );
  DFFR_X1 regBoiz_regfile_reg_2__30_ ( .D(n4458), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__30_) );
  DFFR_X1 regBoiz_regfile_reg_1__30_ ( .D(n4457), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__30_) );
  DFFR_X1 regBoiz_regfile_reg_0__30_ ( .D(n4456), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__30_) );
  DFFR_X1 memBoi_memReg_8__regBoi_curData_reg ( .D(n4455), .CK(clk), .RN(n6873), .Q(wbBusWh[2]), .QN(n5682) );
  DFFR_X1 regBoiz_regfile_reg_31__29_ ( .D(n4454), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__29_) );
  DFFR_X1 regBoiz_regfile_reg_29__29_ ( .D(n4452), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__29_) );
  DFFR_X1 regBoiz_regfile_reg_28__29_ ( .D(n4451), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__29_) );
  DFFR_X1 regBoiz_regfile_reg_27__29_ ( .D(n4450), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__29_) );
  DFFR_X1 regBoiz_regfile_reg_25__29_ ( .D(n4448), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__29_) );
  DFFR_X1 regBoiz_regfile_reg_24__29_ ( .D(n4447), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__29_) );
  DFFR_X1 regBoiz_regfile_reg_23__29_ ( .D(n4446), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__29_) );
  DFFR_X1 regBoiz_regfile_reg_22__29_ ( .D(n4445), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__29_) );
  DFFR_X1 regBoiz_regfile_reg_21__29_ ( .D(n4444), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__29_) );
  DFFR_X1 regBoiz_regfile_reg_20__29_ ( .D(n4443), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__29_) );
  DFFR_X1 regBoiz_regfile_reg_19__29_ ( .D(n4442), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__29_) );
  DFFR_X1 regBoiz_regfile_reg_18__29_ ( .D(n4441), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__29_) );
  DFFR_X1 regBoiz_regfile_reg_17__29_ ( .D(n4440), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__29_) );
  DFFR_X1 regBoiz_regfile_reg_16__29_ ( .D(n4439), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__29_) );
  DFFR_X1 regBoiz_regfile_reg_15__29_ ( .D(n4438), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__29_) );
  DFFR_X1 regBoiz_regfile_reg_13__29_ ( .D(n4436), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__29_) );
  DFFR_X1 regBoiz_regfile_reg_12__29_ ( .D(n4435), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__29_) );
  DFFR_X1 regBoiz_regfile_reg_10__29_ ( .D(n4433), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__29_) );
  DFFR_X1 regBoiz_regfile_reg_9__29_ ( .D(n4432), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_9__29_) );
  DFFR_X1 regBoiz_regfile_reg_8__29_ ( .D(n4431), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__29_) );
  DFFR_X1 regBoiz_regfile_reg_7__29_ ( .D(n4430), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__29_) );
  DFFR_X1 regBoiz_regfile_reg_5__29_ ( .D(n4428), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__29_) );
  DFFR_X1 regBoiz_regfile_reg_4__29_ ( .D(n4427), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__29_) );
  DFFR_X1 regBoiz_regfile_reg_3__29_ ( .D(n4426), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__29_) );
  DFFR_X1 regBoiz_regfile_reg_2__29_ ( .D(n4425), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__29_) );
  DFFR_X1 regBoiz_regfile_reg_1__29_ ( .D(n4424), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__29_) );
  DFFR_X1 regBoiz_regfile_reg_0__29_ ( .D(n4423), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__29_) );
  DFFR_X1 memBoi_memReg_9__regBoi_curData_reg ( .D(n4422), .CK(clk), .RN(n6901), .Q(wbBusWh[3]), .QN(n5668) );
  DFFR_X1 regBoiz_regfile_reg_31__28_ ( .D(n4421), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__28_) );
  DFFR_X1 regBoiz_regfile_reg_30__28_ ( .D(n4420), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__28_) );
  DFFR_X1 regBoiz_regfile_reg_29__28_ ( .D(n4419), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__28_) );
  DFFR_X1 regBoiz_regfile_reg_28__28_ ( .D(n4418), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__28_) );
  DFFR_X1 regBoiz_regfile_reg_27__28_ ( .D(n4417), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__28_) );
  DFFR_X1 regBoiz_regfile_reg_25__28_ ( .D(n4415), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__28_) );
  DFFR_X1 regBoiz_regfile_reg_23__28_ ( .D(n4413), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__28_) );
  DFFR_X1 regBoiz_regfile_reg_21__28_ ( .D(n4411), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__28_) );
  DFFR_X1 regBoiz_regfile_reg_20__28_ ( .D(n4410), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__28_) );
  DFFR_X1 regBoiz_regfile_reg_16__28_ ( .D(n4406), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__28_) );
  DFFR_X1 regBoiz_regfile_reg_15__28_ ( .D(n4405), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__28_) );
  DFFR_X1 regBoiz_regfile_reg_14__28_ ( .D(n4404), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__28_) );
  DFFR_X1 regBoiz_regfile_reg_13__28_ ( .D(n4403), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__28_) );
  DFFR_X1 regBoiz_regfile_reg_12__28_ ( .D(n4402), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__28_) );
  DFFR_X1 regBoiz_regfile_reg_11__28_ ( .D(n4401), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__28_) );
  DFFR_X1 regBoiz_regfile_reg_9__28_ ( .D(n4399), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_9__28_) );
  DFFR_X1 regBoiz_regfile_reg_8__28_ ( .D(n4398), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_8__28_) );
  DFFR_X1 regBoiz_regfile_reg_7__28_ ( .D(n4397), .CK(clk), .RN(n6887), .Q(
        regBoiz_regfile_7__28_) );
  DFFR_X1 regBoiz_regfile_reg_6__28_ ( .D(n4396), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__28_) );
  DFFR_X1 regBoiz_regfile_reg_5__28_ ( .D(n4395), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__28_) );
  DFFR_X1 regBoiz_regfile_reg_4__28_ ( .D(n4394), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__28_) );
  DFFR_X1 regBoiz_regfile_reg_3__28_ ( .D(n4393), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__28_) );
  DFFR_X1 regBoiz_regfile_reg_2__28_ ( .D(n4392), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__28_) );
  DFFR_X1 regBoiz_regfile_reg_1__28_ ( .D(n4391), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__28_) );
  DFFR_X1 regBoiz_regfile_reg_0__28_ ( .D(n4390), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__28_) );
  DFFR_X1 memBoi_memReg_10__regBoi_curData_reg ( .D(n4389), .CK(clk), .RN(
        n6900), .Q(wbBusWh[4]), .QN(n5667) );
  DFFR_X1 regBoiz_regfile_reg_31__27_ ( .D(n4388), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__27_) );
  DFFR_X1 regBoiz_regfile_reg_30__27_ ( .D(n4387), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__27_) );
  DFFR_X1 regBoiz_regfile_reg_29__27_ ( .D(n4386), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__27_) );
  DFFR_X1 regBoiz_regfile_reg_28__27_ ( .D(n4385), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__27_) );
  DFFR_X1 regBoiz_regfile_reg_27__27_ ( .D(n4384), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__27_) );
  DFFR_X1 regBoiz_regfile_reg_26__27_ ( .D(n4383), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__27_), .QN(n5419) );
  DFFR_X1 regBoiz_regfile_reg_25__27_ ( .D(n4382), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__27_) );
  DFFR_X1 regBoiz_regfile_reg_23__27_ ( .D(n4380), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__27_) );
  DFFR_X1 regBoiz_regfile_reg_22__27_ ( .D(n4379), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__27_) );
  DFFR_X1 regBoiz_regfile_reg_21__27_ ( .D(n4378), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__27_) );
  DFFR_X1 regBoiz_regfile_reg_20__27_ ( .D(n4377), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__27_) );
  DFFR_X1 regBoiz_regfile_reg_19__27_ ( .D(n4376), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__27_) );
  DFFR_X1 regBoiz_regfile_reg_18__27_ ( .D(n4375), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__27_), .QN(n5336) );
  DFFR_X1 regBoiz_regfile_reg_17__27_ ( .D(n4374), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__27_) );
  DFFR_X1 regBoiz_regfile_reg_15__27_ ( .D(n4372), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__27_), .QN(n5426) );
  DFFR_X1 regBoiz_regfile_reg_13__27_ ( .D(n4370), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__27_), .QN(n5425) );
  DFFR_X1 regBoiz_regfile_reg_12__27_ ( .D(n4369), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__27_) );
  DFFR_X1 regBoiz_regfile_reg_11__27_ ( .D(n4368), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__27_), .QN(n5424) );
  DFFR_X1 regBoiz_regfile_reg_9__27_ ( .D(n4366), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_9__27_), .QN(n5423) );
  DFFR_X1 regBoiz_regfile_reg_8__27_ ( .D(n4365), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__27_) );
  DFFR_X1 regBoiz_regfile_reg_7__27_ ( .D(n4364), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__27_), .QN(n5340) );
  DFFR_X1 regBoiz_regfile_reg_6__27_ ( .D(n4363), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__27_) );
  DFFR_X1 regBoiz_regfile_reg_5__27_ ( .D(n4362), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__27_), .QN(n5339) );
  DFFR_X1 regBoiz_regfile_reg_4__27_ ( .D(n4361), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__27_) );
  DFFR_X1 regBoiz_regfile_reg_3__27_ ( .D(n4360), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__27_), .QN(n5338) );
  DFFR_X1 regBoiz_regfile_reg_2__27_ ( .D(n4359), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__27_) );
  DFFR_X1 regBoiz_regfile_reg_1__27_ ( .D(n4358), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__27_), .QN(n5337) );
  DFFR_X1 regBoiz_regfile_reg_0__27_ ( .D(n4357), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__27_) );
  DFFR_X1 memBoi_memReg_11__regBoi_curData_reg ( .D(n4356), .CK(clk), .RN(
        n6875), .Q(wbBusWh[5]), .QN(n5666) );
  DFFR_X1 regBoiz_regfile_reg_31__26_ ( .D(n4355), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__26_) );
  DFFR_X1 regBoiz_regfile_reg_30__26_ ( .D(n4354), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__26_) );
  DFFR_X1 regBoiz_regfile_reg_29__26_ ( .D(n4353), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__26_) );
  DFFR_X1 regBoiz_regfile_reg_28__26_ ( .D(n4352), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__26_) );
  DFFR_X1 regBoiz_regfile_reg_27__26_ ( .D(n4351), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__26_) );
  DFFR_X1 regBoiz_regfile_reg_26__26_ ( .D(n4350), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__26_) );
  DFFR_X1 regBoiz_regfile_reg_25__26_ ( .D(n4349), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__26_) );
  DFFR_X1 regBoiz_regfile_reg_24__26_ ( .D(n4348), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__26_) );
  DFFR_X1 regBoiz_regfile_reg_23__26_ ( .D(n4347), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__26_) );
  DFFR_X1 regBoiz_regfile_reg_22__26_ ( .D(n4346), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__26_) );
  DFFR_X1 regBoiz_regfile_reg_21__26_ ( .D(n4345), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__26_) );
  DFFR_X1 regBoiz_regfile_reg_20__26_ ( .D(n4344), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__26_) );
  DFFR_X1 regBoiz_regfile_reg_19__26_ ( .D(n4343), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__26_) );
  DFFR_X1 regBoiz_regfile_reg_18__26_ ( .D(n4342), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__26_) );
  DFFR_X1 regBoiz_regfile_reg_17__26_ ( .D(n4341), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__26_) );
  DFFR_X1 regBoiz_regfile_reg_16__26_ ( .D(n4340), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__26_) );
  DFFR_X1 regBoiz_regfile_reg_14__26_ ( .D(n4338), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__26_) );
  DFFR_X1 regBoiz_regfile_reg_13__26_ ( .D(n4337), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__26_), .QN(n5588) );
  DFFR_X1 regBoiz_regfile_reg_12__26_ ( .D(n4336), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__26_) );
  DFFR_X1 regBoiz_regfile_reg_11__26_ ( .D(n4335), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__26_), .QN(n5341) );
  DFFR_X1 regBoiz_regfile_reg_10__26_ ( .D(n4334), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__26_), .QN(n6141) );
  DFFR_X1 regBoiz_regfile_reg_9__26_ ( .D(n4333), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_9__26_), .QN(n5589) );
  DFFR_X1 regBoiz_regfile_reg_8__26_ ( .D(n4332), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_8__26_) );
  DFFR_X1 regBoiz_regfile_reg_7__26_ ( .D(n4331), .CK(clk), .RN(n6900), .Q(
        regBoiz_regfile_7__26_), .QN(n5931) );
  DFFR_X1 regBoiz_regfile_reg_6__26_ ( .D(n4330), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__26_) );
  DFFR_X1 regBoiz_regfile_reg_5__26_ ( .D(n4329), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__26_), .QN(n5382) );
  DFFR_X1 regBoiz_regfile_reg_4__26_ ( .D(n4328), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__26_) );
  DFFR_X1 regBoiz_regfile_reg_3__26_ ( .D(n4327), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__26_), .QN(n5578) );
  DFFR_X1 regBoiz_regfile_reg_2__26_ ( .D(n4326), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__26_), .QN(n6142) );
  DFFR_X1 regBoiz_regfile_reg_1__26_ ( .D(n4325), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__26_), .QN(n5383) );
  DFFR_X1 regBoiz_regfile_reg_0__26_ ( .D(n4324), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__26_) );
  DFFR_X1 memBoi_memReg_12__regBoi_curData_reg ( .D(n4323), .CK(clk), .RN(
        n6900), .Q(wbBusWh[6]), .QN(n5665) );
  DFFR_X1 regBoiz_regfile_reg_31__25_ ( .D(n4322), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__25_) );
  DFFR_X1 regBoiz_regfile_reg_30__25_ ( .D(n4321), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__25_) );
  DFFR_X1 regBoiz_regfile_reg_29__25_ ( .D(n4320), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__25_) );
  DFFR_X1 regBoiz_regfile_reg_28__25_ ( .D(n4319), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__25_) );
  DFFR_X1 regBoiz_regfile_reg_27__25_ ( .D(n4318), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__25_) );
  DFFR_X1 regBoiz_regfile_reg_26__25_ ( .D(n4317), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__25_) );
  DFFR_X1 regBoiz_regfile_reg_25__25_ ( .D(n4316), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__25_) );
  DFFR_X1 regBoiz_regfile_reg_24__25_ ( .D(n4315), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__25_) );
  DFFR_X1 regBoiz_regfile_reg_23__25_ ( .D(n4314), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__25_) );
  DFFR_X1 regBoiz_regfile_reg_22__25_ ( .D(n4313), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__25_) );
  DFFR_X1 regBoiz_regfile_reg_21__25_ ( .D(n4312), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__25_) );
  DFFR_X1 regBoiz_regfile_reg_20__25_ ( .D(n4311), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__25_) );
  DFFR_X1 regBoiz_regfile_reg_19__25_ ( .D(n4310), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__25_) );
  DFFR_X1 regBoiz_regfile_reg_18__25_ ( .D(n4309), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__25_) );
  DFFR_X1 regBoiz_regfile_reg_17__25_ ( .D(n4308), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__25_) );
  DFFR_X1 regBoiz_regfile_reg_16__25_ ( .D(n4307), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__25_) );
  DFFR_X1 regBoiz_regfile_reg_15__25_ ( .D(n4306), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__25_) );
  DFFR_X1 regBoiz_regfile_reg_14__25_ ( .D(n4305), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__25_) );
  DFFR_X1 regBoiz_regfile_reg_13__25_ ( .D(n4304), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__25_) );
  DFFR_X1 regBoiz_regfile_reg_12__25_ ( .D(n4303), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__25_) );
  DFFR_X1 regBoiz_regfile_reg_11__25_ ( .D(n4302), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__25_) );
  DFFR_X1 regBoiz_regfile_reg_10__25_ ( .D(n4301), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__25_) );
  DFFR_X1 regBoiz_regfile_reg_9__25_ ( .D(n4300), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_9__25_) );
  DFFR_X1 regBoiz_regfile_reg_8__25_ ( .D(n4299), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__25_) );
  DFFR_X1 regBoiz_regfile_reg_7__25_ ( .D(n4298), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__25_) );
  DFFR_X1 regBoiz_regfile_reg_6__25_ ( .D(n4297), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__25_) );
  DFFR_X1 regBoiz_regfile_reg_5__25_ ( .D(n4296), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__25_) );
  DFFR_X1 regBoiz_regfile_reg_4__25_ ( .D(n4295), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__25_) );
  DFFR_X1 regBoiz_regfile_reg_3__25_ ( .D(n4294), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__25_) );
  DFFR_X1 regBoiz_regfile_reg_2__25_ ( .D(n4293), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__25_) );
  DFFR_X1 regBoiz_regfile_reg_1__25_ ( .D(n4292), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__25_) );
  DFFR_X1 regBoiz_regfile_reg_0__25_ ( .D(n4291), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__25_) );
  DFFR_X1 memBoi_memReg_13__regBoi_curData_reg ( .D(n13677), .CK(clk), .RN(
        n6875), .Q(wbBusWh[7]), .QN(n5664) );
  DFFR_X1 regBoiz_regfile_reg_31__24_ ( .D(n4289), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__24_) );
  DFFR_X1 regBoiz_regfile_reg_30__24_ ( .D(n4288), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__24_) );
  DFFR_X1 regBoiz_regfile_reg_29__24_ ( .D(n4287), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__24_) );
  DFFR_X1 regBoiz_regfile_reg_28__24_ ( .D(n4286), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__24_) );
  DFFR_X1 regBoiz_regfile_reg_27__24_ ( .D(n4285), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__24_) );
  DFFR_X1 regBoiz_regfile_reg_26__24_ ( .D(n4284), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__24_) );
  DFFR_X1 regBoiz_regfile_reg_25__24_ ( .D(n4283), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__24_) );
  DFFR_X1 regBoiz_regfile_reg_24__24_ ( .D(n4282), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__24_) );
  DFFR_X1 regBoiz_regfile_reg_23__24_ ( .D(n4281), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__24_) );
  DFFR_X1 regBoiz_regfile_reg_22__24_ ( .D(n4280), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__24_) );
  DFFR_X1 regBoiz_regfile_reg_21__24_ ( .D(n4279), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__24_) );
  DFFR_X1 regBoiz_regfile_reg_20__24_ ( .D(n4278), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__24_) );
  DFFR_X1 regBoiz_regfile_reg_19__24_ ( .D(n4277), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__24_) );
  DFFR_X1 regBoiz_regfile_reg_18__24_ ( .D(n4276), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__24_) );
  DFFR_X1 regBoiz_regfile_reg_17__24_ ( .D(n4275), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__24_) );
  DFFR_X1 regBoiz_regfile_reg_16__24_ ( .D(n4274), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__24_) );
  DFFR_X1 regBoiz_regfile_reg_15__24_ ( .D(n4273), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__24_) );
  DFFR_X1 regBoiz_regfile_reg_14__24_ ( .D(n4272), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__24_) );
  DFFR_X1 regBoiz_regfile_reg_13__24_ ( .D(n4271), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__24_) );
  DFFR_X1 regBoiz_regfile_reg_12__24_ ( .D(n4270), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__24_) );
  DFFR_X1 regBoiz_regfile_reg_11__24_ ( .D(n4269), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__24_) );
  DFFR_X1 regBoiz_regfile_reg_10__24_ ( .D(n4268), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__24_) );
  DFFR_X1 regBoiz_regfile_reg_9__24_ ( .D(n4267), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_9__24_) );
  DFFR_X1 regBoiz_regfile_reg_8__24_ ( .D(n4266), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_8__24_) );
  DFFR_X1 regBoiz_regfile_reg_7__24_ ( .D(n4265), .CK(clk), .RN(n6901), .Q(
        regBoiz_regfile_7__24_) );
  DFFR_X1 regBoiz_regfile_reg_6__24_ ( .D(n4264), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__24_) );
  DFFR_X1 regBoiz_regfile_reg_5__24_ ( .D(n4263), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__24_) );
  DFFR_X1 regBoiz_regfile_reg_4__24_ ( .D(n4262), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__24_) );
  DFFR_X1 regBoiz_regfile_reg_3__24_ ( .D(n4261), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__24_) );
  DFFR_X1 regBoiz_regfile_reg_2__24_ ( .D(n4260), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__24_) );
  DFFR_X1 regBoiz_regfile_reg_1__24_ ( .D(n4259), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__24_) );
  DFFR_X1 regBoiz_regfile_reg_0__24_ ( .D(n4258), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__24_) );
  DFFR_X1 memBoi_memReg_14__regBoi_curData_reg ( .D(n4257), .CK(clk), .RN(
        n6900), .Q(wbBusWh[8]), .QN(n5663) );
  DFFR_X1 regBoiz_regfile_reg_29__23_ ( .D(n4254), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__23_), .QN(n6190) );
  DFFR_X1 regBoiz_regfile_reg_28__23_ ( .D(n4253), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__23_), .QN(n6369) );
  DFFR_X1 regBoiz_regfile_reg_25__23_ ( .D(n4250), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__23_), .QN(n6189) );
  DFFR_X1 regBoiz_regfile_reg_21__23_ ( .D(n4246), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__23_) );
  DFFR_X1 regBoiz_regfile_reg_20__23_ ( .D(n4245), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__23_), .QN(n6368) );
  DFFR_X1 regBoiz_regfile_reg_19__23_ ( .D(n4244), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__23_) );
  DFFR_X1 regBoiz_regfile_reg_17__23_ ( .D(n4242), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__23_) );
  DFFR_X1 regBoiz_regfile_reg_16__23_ ( .D(n4241), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__23_) );
  DFFR_X1 regBoiz_regfile_reg_14__23_ ( .D(n4239), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__23_) );
  DFFR_X1 regBoiz_regfile_reg_13__23_ ( .D(n4238), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__23_) );
  DFFR_X1 regBoiz_regfile_reg_12__23_ ( .D(n4237), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__23_) );
  DFFR_X1 regBoiz_regfile_reg_11__23_ ( .D(n4236), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__23_) );
  DFFR_X1 regBoiz_regfile_reg_10__23_ ( .D(n4235), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__23_) );
  DFFR_X1 regBoiz_regfile_reg_9__23_ ( .D(n4234), .CK(clk), .RN(n6891), .Q(
        regBoiz_regfile_9__23_) );
  DFFR_X1 regBoiz_regfile_reg_8__23_ ( .D(n4233), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__23_) );
  DFFR_X1 regBoiz_regfile_reg_7__23_ ( .D(n4232), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__23_) );
  DFFR_X1 regBoiz_regfile_reg_6__23_ ( .D(n4231), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__23_) );
  DFFR_X1 regBoiz_regfile_reg_5__23_ ( .D(n4230), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__23_) );
  DFFR_X1 regBoiz_regfile_reg_4__23_ ( .D(n4229), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__23_) );
  DFFR_X1 regBoiz_regfile_reg_3__23_ ( .D(n4228), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__23_) );
  DFFR_X1 regBoiz_regfile_reg_2__23_ ( .D(n4227), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__23_) );
  DFFR_X1 regBoiz_regfile_reg_1__23_ ( .D(n4226), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__23_) );
  DFFR_X1 regBoiz_regfile_reg_0__23_ ( .D(n4225), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__23_) );
  DFFR_X1 memBoi_memReg_15__regBoi_curData_reg ( .D(n4224), .CK(clk), .RN(
        n6874), .Q(wbBusWh[9]), .QN(n5662) );
  DFFR_X1 regBoiz_regfile_reg_31__22_ ( .D(n4223), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__22_) );
  DFFR_X1 regBoiz_regfile_reg_30__22_ ( .D(n4222), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__22_) );
  DFFR_X1 regBoiz_regfile_reg_29__22_ ( .D(n4221), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_29__22_) );
  DFFR_X1 regBoiz_regfile_reg_28__22_ ( .D(n4220), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__22_) );
  DFFR_X1 regBoiz_regfile_reg_27__22_ ( .D(n4219), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__22_) );
  DFFR_X1 regBoiz_regfile_reg_26__22_ ( .D(n4218), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__22_) );
  DFFR_X1 regBoiz_regfile_reg_25__22_ ( .D(n4217), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__22_) );
  DFFR_X1 regBoiz_regfile_reg_24__22_ ( .D(n4216), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__22_) );
  DFFR_X1 regBoiz_regfile_reg_23__22_ ( .D(n4215), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__22_) );
  DFFR_X1 regBoiz_regfile_reg_22__22_ ( .D(n4214), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__22_) );
  DFFR_X1 regBoiz_regfile_reg_21__22_ ( .D(n4213), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__22_) );
  DFFR_X1 regBoiz_regfile_reg_20__22_ ( .D(n4212), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__22_) );
  DFFR_X1 regBoiz_regfile_reg_19__22_ ( .D(n4211), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__22_) );
  DFFR_X1 regBoiz_regfile_reg_18__22_ ( .D(n4210), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__22_) );
  DFFR_X1 regBoiz_regfile_reg_17__22_ ( .D(n4209), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__22_) );
  DFFR_X1 regBoiz_regfile_reg_16__22_ ( .D(n4208), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__22_) );
  DFFR_X1 regBoiz_regfile_reg_14__22_ ( .D(n4206), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__22_) );
  DFFR_X1 regBoiz_regfile_reg_13__22_ ( .D(n4205), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__22_) );
  DFFR_X1 regBoiz_regfile_reg_12__22_ ( .D(n4204), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__22_) );
  DFFR_X1 regBoiz_regfile_reg_11__22_ ( .D(n4203), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__22_) );
  DFFR_X1 regBoiz_regfile_reg_10__22_ ( .D(n4202), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__22_) );
  DFFR_X1 regBoiz_regfile_reg_9__22_ ( .D(n4201), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_9__22_) );
  DFFR_X1 regBoiz_regfile_reg_8__22_ ( .D(n4200), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_8__22_) );
  DFFR_X1 regBoiz_regfile_reg_7__22_ ( .D(n4199), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_7__22_) );
  DFFR_X1 regBoiz_regfile_reg_6__22_ ( .D(n4198), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__22_) );
  DFFR_X1 regBoiz_regfile_reg_5__22_ ( .D(n4197), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__22_) );
  DFFR_X1 regBoiz_regfile_reg_4__22_ ( .D(n4196), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__22_) );
  DFFR_X1 regBoiz_regfile_reg_3__22_ ( .D(n4195), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__22_) );
  DFFR_X1 regBoiz_regfile_reg_2__22_ ( .D(n4194), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__22_) );
  DFFR_X1 regBoiz_regfile_reg_1__22_ ( .D(n4193), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__22_) );
  DFFR_X1 regBoiz_regfile_reg_0__22_ ( .D(n4192), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__22_) );
  DFFR_X1 memBoi_memReg_16__regBoi_curData_reg ( .D(n4191), .CK(clk), .RN(
        n6900), .Q(wbBusWh[10]), .QN(n5661) );
  DFFR_X1 regBoiz_regfile_reg_31__21_ ( .D(n4190), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__21_) );
  DFFR_X1 regBoiz_regfile_reg_30__21_ ( .D(n4189), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__21_) );
  DFFR_X1 regBoiz_regfile_reg_29__21_ ( .D(n4188), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__21_) );
  DFFR_X1 regBoiz_regfile_reg_28__21_ ( .D(n4187), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__21_) );
  DFFR_X1 regBoiz_regfile_reg_27__21_ ( .D(n4186), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__21_), .QN(n5549) );
  DFFR_X1 regBoiz_regfile_reg_25__21_ ( .D(n4184), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__21_), .QN(n5547) );
  DFFR_X1 regBoiz_regfile_reg_23__21_ ( .D(n4182), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__21_) );
  DFFR_X1 regBoiz_regfile_reg_22__21_ ( .D(n4181), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__21_) );
  DFFR_X1 regBoiz_regfile_reg_21__21_ ( .D(n4180), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__21_) );
  DFFR_X1 regBoiz_regfile_reg_20__21_ ( .D(n4179), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__21_) );
  DFFR_X1 regBoiz_regfile_reg_15__21_ ( .D(n4174), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__21_) );
  DFFR_X1 regBoiz_regfile_reg_14__21_ ( .D(n4173), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__21_) );
  DFFR_X1 regBoiz_regfile_reg_13__21_ ( .D(n4172), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__21_) );
  DFFR_X1 regBoiz_regfile_reg_12__21_ ( .D(n4171), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__21_) );
  DFFR_X1 regBoiz_regfile_reg_11__21_ ( .D(n4170), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__21_), .QN(n5548) );
  DFFR_X1 regBoiz_regfile_reg_10__21_ ( .D(n4169), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__21_), .QN(n5532) );
  DFFR_X1 regBoiz_regfile_reg_9__21_ ( .D(n4168), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_9__21_), .QN(n5546) );
  DFFR_X1 regBoiz_regfile_reg_7__21_ ( .D(n4166), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__21_) );
  DFFR_X1 regBoiz_regfile_reg_6__21_ ( .D(n4165), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__21_) );
  DFFR_X1 regBoiz_regfile_reg_5__21_ ( .D(n4164), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__21_) );
  DFFR_X1 regBoiz_regfile_reg_4__21_ ( .D(n4163), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__21_) );
  DFFR_X1 regBoiz_regfile_reg_3__21_ ( .D(n4162), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__21_), .QN(n5550) );
  DFFR_X1 regBoiz_regfile_reg_2__21_ ( .D(n4161), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__21_), .QN(n5533) );
  DFFR_X1 regBoiz_regfile_reg_1__21_ ( .D(n4160), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__21_), .QN(n5637) );
  DFFR_X1 memBoi_memReg_17__regBoi_curData_reg ( .D(n4158), .CK(clk), .RN(
        n6874), .Q(wbBusWh[11]), .QN(n5660) );
  DFFR_X1 regBoiz_regfile_reg_31__20_ ( .D(n4157), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__20_) );
  DFFR_X1 regBoiz_regfile_reg_29__20_ ( .D(n4155), .CK(clk), .RN(n6898), .Q(
        regBoiz_regfile_29__20_) );
  DFFR_X1 regBoiz_regfile_reg_28__20_ ( .D(n4154), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__20_) );
  DFFR_X1 regBoiz_regfile_reg_27__20_ ( .D(n4153), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__20_) );
  DFFR_X1 regBoiz_regfile_reg_26__20_ ( .D(n4152), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__20_) );
  DFFR_X1 regBoiz_regfile_reg_25__20_ ( .D(n4151), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__20_) );
  DFFR_X1 regBoiz_regfile_reg_24__20_ ( .D(n4150), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__20_) );
  DFFR_X1 regBoiz_regfile_reg_23__20_ ( .D(n4149), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__20_) );
  DFFR_X1 regBoiz_regfile_reg_22__20_ ( .D(n4148), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__20_) );
  DFFR_X1 regBoiz_regfile_reg_21__20_ ( .D(n4147), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__20_) );
  DFFR_X1 regBoiz_regfile_reg_20__20_ ( .D(n4146), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__20_) );
  DFFR_X1 regBoiz_regfile_reg_19__20_ ( .D(n4145), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__20_) );
  DFFR_X1 regBoiz_regfile_reg_18__20_ ( .D(n4144), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__20_) );
  DFFR_X1 regBoiz_regfile_reg_17__20_ ( .D(n4143), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__20_) );
  DFFR_X1 regBoiz_regfile_reg_16__20_ ( .D(n4142), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__20_) );
  DFFR_X1 regBoiz_regfile_reg_15__20_ ( .D(n4141), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__20_) );
  DFFR_X1 regBoiz_regfile_reg_14__20_ ( .D(n4140), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__20_) );
  DFFR_X1 regBoiz_regfile_reg_13__20_ ( .D(n4139), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__20_) );
  DFFR_X1 regBoiz_regfile_reg_12__20_ ( .D(n4138), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__20_) );
  DFFR_X1 regBoiz_regfile_reg_11__20_ ( .D(n4137), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__20_) );
  DFFR_X1 regBoiz_regfile_reg_10__20_ ( .D(n4136), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__20_) );
  DFFR_X1 regBoiz_regfile_reg_9__20_ ( .D(n4135), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_9__20_) );
  DFFR_X1 regBoiz_regfile_reg_8__20_ ( .D(n4134), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_8__20_) );
  DFFR_X1 regBoiz_regfile_reg_7__20_ ( .D(n4133), .CK(clk), .RN(n6888), .Q(
        regBoiz_regfile_7__20_) );
  DFFR_X1 regBoiz_regfile_reg_6__20_ ( .D(n4132), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__20_) );
  DFFR_X1 regBoiz_regfile_reg_5__20_ ( .D(n4131), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__20_) );
  DFFR_X1 regBoiz_regfile_reg_4__20_ ( .D(n4130), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__20_) );
  DFFR_X1 regBoiz_regfile_reg_3__20_ ( .D(n4129), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__20_) );
  DFFR_X1 regBoiz_regfile_reg_2__20_ ( .D(n4128), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__20_) );
  DFFR_X1 regBoiz_regfile_reg_1__20_ ( .D(n4127), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__20_) );
  DFFR_X1 regBoiz_regfile_reg_0__20_ ( .D(n4126), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__20_) );
  DFFR_X1 memBoi_memReg_18__regBoi_curData_reg ( .D(n4125), .CK(clk), .RN(
        n6900), .Q(wbBusWh[12]), .QN(n5658) );
  DFFR_X1 regBoiz_regfile_reg_31__19_ ( .D(n4124), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__19_) );
  DFFR_X1 regBoiz_regfile_reg_30__19_ ( .D(n4123), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__19_) );
  DFFR_X1 regBoiz_regfile_reg_29__19_ ( .D(n4122), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_29__19_) );
  DFFR_X1 regBoiz_regfile_reg_28__19_ ( .D(n4121), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__19_) );
  DFFR_X1 regBoiz_regfile_reg_27__19_ ( .D(n4120), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__19_) );
  DFFR_X1 regBoiz_regfile_reg_26__19_ ( .D(n4119), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__19_), .QN(n5567) );
  DFFR_X1 regBoiz_regfile_reg_25__19_ ( .D(n4118), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__19_) );
  DFFR_X1 regBoiz_regfile_reg_24__19_ ( .D(n4117), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__19_) );
  DFFR_X1 regBoiz_regfile_reg_23__19_ ( .D(n4116), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__19_) );
  DFFR_X1 regBoiz_regfile_reg_22__19_ ( .D(n4115), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__19_) );
  DFFR_X1 regBoiz_regfile_reg_21__19_ ( .D(n4114), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__19_) );
  DFFR_X1 regBoiz_regfile_reg_20__19_ ( .D(n4113), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__19_) );
  DFFR_X1 regBoiz_regfile_reg_19__19_ ( .D(n4112), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__19_) );
  DFFR_X1 regBoiz_regfile_reg_18__19_ ( .D(n4111), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__19_), .QN(n5566) );
  DFFR_X1 regBoiz_regfile_reg_17__19_ ( .D(n4110), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__19_) );
  DFFR_X1 regBoiz_regfile_reg_16__19_ ( .D(n4109), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__19_) );
  DFFR_X1 regBoiz_regfile_reg_15__19_ ( .D(n4108), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__19_) );
  DFFR_X1 regBoiz_regfile_reg_14__19_ ( .D(n4107), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__19_) );
  DFFR_X1 regBoiz_regfile_reg_13__19_ ( .D(n4106), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__19_) );
  DFFR_X1 regBoiz_regfile_reg_12__19_ ( .D(n4105), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__19_) );
  DFFR_X1 regBoiz_regfile_reg_11__19_ ( .D(n4104), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__19_) );
  DFFR_X1 regBoiz_regfile_reg_10__19_ ( .D(n4103), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__19_) );
  DFFR_X1 regBoiz_regfile_reg_9__19_ ( .D(n4102), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_9__19_) );
  DFFR_X1 regBoiz_regfile_reg_8__19_ ( .D(n4101), .CK(clk), .RN(n6886), .Q(
        regBoiz_regfile_8__19_), .QN(n5568) );
  DFFR_X1 regBoiz_regfile_reg_7__19_ ( .D(n4100), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_7__19_) );
  DFFR_X1 regBoiz_regfile_reg_6__19_ ( .D(n4099), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__19_) );
  DFFR_X1 regBoiz_regfile_reg_5__19_ ( .D(n4098), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__19_) );
  DFFR_X1 regBoiz_regfile_reg_4__19_ ( .D(n4097), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__19_) );
  DFFR_X1 regBoiz_regfile_reg_3__19_ ( .D(n4096), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__19_) );
  DFFR_X1 regBoiz_regfile_reg_2__19_ ( .D(n4095), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__19_) );
  DFFR_X1 regBoiz_regfile_reg_1__19_ ( .D(n4094), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__19_) );
  DFFR_X1 regBoiz_regfile_reg_0__19_ ( .D(n4093), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__19_), .QN(n5582) );
  DFFR_X1 memBoi_memReg_19__regBoi_curData_reg ( .D(n4092), .CK(clk), .RN(
        n6874), .Q(wbBusWh[13]), .QN(n5657) );
  DFFR_X1 regBoiz_regfile_reg_31__18_ ( .D(n4091), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__18_) );
  DFFR_X1 regBoiz_regfile_reg_30__18_ ( .D(n4090), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__18_) );
  DFFR_X1 regBoiz_regfile_reg_29__18_ ( .D(n4089), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__18_) );
  DFFR_X1 regBoiz_regfile_reg_28__18_ ( .D(n4088), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__18_) );
  DFFR_X1 regBoiz_regfile_reg_27__18_ ( .D(n4087), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__18_) );
  DFFR_X1 regBoiz_regfile_reg_26__18_ ( .D(n4086), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__18_) );
  DFFR_X1 regBoiz_regfile_reg_25__18_ ( .D(n4085), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__18_) );
  DFFR_X1 regBoiz_regfile_reg_23__18_ ( .D(n4083), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__18_) );
  DFFR_X1 regBoiz_regfile_reg_22__18_ ( .D(n4082), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__18_) );
  DFFR_X1 regBoiz_regfile_reg_21__18_ ( .D(n4081), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__18_) );
  DFFR_X1 regBoiz_regfile_reg_20__18_ ( .D(n4080), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__18_) );
  DFFR_X1 regBoiz_regfile_reg_19__18_ ( .D(n4079), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__18_) );
  DFFR_X1 regBoiz_regfile_reg_18__18_ ( .D(n4078), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__18_) );
  DFFR_X1 regBoiz_regfile_reg_17__18_ ( .D(n4077), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__18_) );
  DFFR_X1 regBoiz_regfile_reg_16__18_ ( .D(n4076), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__18_) );
  DFFR_X1 regBoiz_regfile_reg_15__18_ ( .D(n4075), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__18_) );
  DFFR_X1 regBoiz_regfile_reg_14__18_ ( .D(n4074), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__18_) );
  DFFR_X1 regBoiz_regfile_reg_13__18_ ( .D(n4073), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__18_) );
  DFFR_X1 regBoiz_regfile_reg_12__18_ ( .D(n4072), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__18_) );
  DFFR_X1 regBoiz_regfile_reg_11__18_ ( .D(n4071), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__18_) );
  DFFR_X1 regBoiz_regfile_reg_10__18_ ( .D(n4070), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__18_) );
  DFFR_X1 regBoiz_regfile_reg_9__18_ ( .D(n4069), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_9__18_) );
  DFFR_X1 regBoiz_regfile_reg_8__18_ ( .D(n4068), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__18_) );
  DFFR_X1 regBoiz_regfile_reg_7__18_ ( .D(n4067), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__18_) );
  DFFR_X1 regBoiz_regfile_reg_6__18_ ( .D(n4066), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__18_) );
  DFFR_X1 regBoiz_regfile_reg_5__18_ ( .D(n4065), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__18_) );
  DFFR_X1 regBoiz_regfile_reg_4__18_ ( .D(n4064), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__18_) );
  DFFR_X1 regBoiz_regfile_reg_3__18_ ( .D(n4063), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__18_) );
  DFFR_X1 regBoiz_regfile_reg_2__18_ ( .D(n4062), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__18_) );
  DFFR_X1 regBoiz_regfile_reg_1__18_ ( .D(n4061), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__18_) );
  DFFR_X1 regBoiz_regfile_reg_0__18_ ( .D(n4060), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__18_) );
  DFFR_X1 memBoi_memReg_20__regBoi_curData_reg ( .D(n4059), .CK(clk), .RN(
        n6874), .Q(wbBusWh[14]), .QN(n5656) );
  DFFR_X1 regBoiz_regfile_reg_31__17_ ( .D(n4058), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__17_) );
  DFFR_X1 regBoiz_regfile_reg_30__17_ ( .D(n4057), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__17_) );
  DFFR_X1 regBoiz_regfile_reg_29__17_ ( .D(n4056), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_29__17_) );
  DFFR_X1 regBoiz_regfile_reg_28__17_ ( .D(n4055), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__17_) );
  DFFR_X1 regBoiz_regfile_reg_27__17_ ( .D(n4054), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__17_) );
  DFFR_X1 regBoiz_regfile_reg_26__17_ ( .D(n4053), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__17_) );
  DFFR_X1 regBoiz_regfile_reg_25__17_ ( .D(n4052), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__17_) );
  DFFR_X1 regBoiz_regfile_reg_24__17_ ( .D(n4051), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__17_) );
  DFFR_X1 regBoiz_regfile_reg_23__17_ ( .D(n4050), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__17_) );
  DFFR_X1 regBoiz_regfile_reg_22__17_ ( .D(n4049), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__17_) );
  DFFR_X1 regBoiz_regfile_reg_21__17_ ( .D(n4048), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__17_) );
  DFFR_X1 regBoiz_regfile_reg_20__17_ ( .D(n4047), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__17_) );
  DFFR_X1 regBoiz_regfile_reg_19__17_ ( .D(n4046), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__17_) );
  DFFR_X1 regBoiz_regfile_reg_18__17_ ( .D(n4045), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__17_) );
  DFFR_X1 regBoiz_regfile_reg_17__17_ ( .D(n4044), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__17_) );
  DFFR_X1 regBoiz_regfile_reg_16__17_ ( .D(n4043), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__17_) );
  DFFR_X1 regBoiz_regfile_reg_15__17_ ( .D(n4042), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__17_) );
  DFFR_X1 regBoiz_regfile_reg_14__17_ ( .D(n4041), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__17_) );
  DFFR_X1 regBoiz_regfile_reg_13__17_ ( .D(n4040), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__17_) );
  DFFR_X1 regBoiz_regfile_reg_12__17_ ( .D(n4039), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__17_) );
  DFFR_X1 regBoiz_regfile_reg_11__17_ ( .D(n4038), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__17_) );
  DFFR_X1 regBoiz_regfile_reg_10__17_ ( .D(n4037), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__17_) );
  DFFR_X1 regBoiz_regfile_reg_9__17_ ( .D(n4036), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_9__17_) );
  DFFR_X1 regBoiz_regfile_reg_8__17_ ( .D(n4035), .CK(clk), .RN(n6880), .Q(
        regBoiz_regfile_8__17_) );
  DFFR_X1 regBoiz_regfile_reg_7__17_ ( .D(n4034), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_7__17_) );
  DFFR_X1 regBoiz_regfile_reg_6__17_ ( .D(n4033), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__17_) );
  DFFR_X1 regBoiz_regfile_reg_5__17_ ( .D(n4032), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__17_) );
  DFFR_X1 regBoiz_regfile_reg_4__17_ ( .D(n4031), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__17_) );
  DFFR_X1 regBoiz_regfile_reg_3__17_ ( .D(n4030), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__17_) );
  DFFR_X1 regBoiz_regfile_reg_2__17_ ( .D(n4029), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__17_) );
  DFFR_X1 regBoiz_regfile_reg_1__17_ ( .D(n4028), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__17_) );
  DFFR_X1 regBoiz_regfile_reg_0__17_ ( .D(n4027), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__17_) );
  DFFR_X1 memBoi_memReg_21__regBoi_curData_reg ( .D(n4026), .CK(clk), .RN(
        n6900), .Q(wbBusWh[15]), .QN(n5655) );
  DFFR_X1 regBoiz_regfile_reg_30__16_ ( .D(n4024), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__16_) );
  DFFR_X1 regBoiz_regfile_reg_29__16_ ( .D(n4023), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_29__16_) );
  DFFR_X1 regBoiz_regfile_reg_28__16_ ( .D(n4022), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__16_) );
  DFFR_X1 regBoiz_regfile_reg_27__16_ ( .D(n4021), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__16_) );
  DFFR_X1 regBoiz_regfile_reg_26__16_ ( .D(n4020), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_26__16_) );
  DFFR_X1 regBoiz_regfile_reg_25__16_ ( .D(n4019), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__16_) );
  DFFR_X1 regBoiz_regfile_reg_24__16_ ( .D(n4018), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__16_) );
  DFFR_X1 regBoiz_regfile_reg_23__16_ ( .D(n4017), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_23__16_) );
  DFFR_X1 regBoiz_regfile_reg_22__16_ ( .D(n4016), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__16_) );
  DFFR_X1 regBoiz_regfile_reg_21__16_ ( .D(n4015), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__16_) );
  DFFR_X1 regBoiz_regfile_reg_20__16_ ( .D(n4014), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_20__16_) );
  DFFR_X1 regBoiz_regfile_reg_19__16_ ( .D(n4013), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__16_) );
  DFFR_X1 regBoiz_regfile_reg_18__16_ ( .D(n4012), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_18__16_) );
  DFFR_X1 regBoiz_regfile_reg_17__16_ ( .D(n4011), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__16_) );
  DFFR_X1 regBoiz_regfile_reg_16__16_ ( .D(n4010), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__16_) );
  DFFR_X1 regBoiz_regfile_reg_13__16_ ( .D(n4007), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__16_) );
  DFFR_X1 regBoiz_regfile_reg_12__16_ ( .D(n4006), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_12__16_) );
  DFFR_X1 regBoiz_regfile_reg_11__16_ ( .D(n4005), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__16_) );
  DFFR_X1 regBoiz_regfile_reg_10__16_ ( .D(n4004), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__16_) );
  DFFR_X1 regBoiz_regfile_reg_9__16_ ( .D(n4003), .CK(clk), .RN(n6892), .Q(
        regBoiz_regfile_9__16_) );
  DFFR_X1 regBoiz_regfile_reg_8__16_ ( .D(n4002), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_8__16_) );
  DFFR_X1 regBoiz_regfile_reg_7__16_ ( .D(n4001), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__16_) );
  DFFR_X1 regBoiz_regfile_reg_6__16_ ( .D(n4000), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__16_) );
  DFFR_X1 regBoiz_regfile_reg_5__16_ ( .D(n3999), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_5__16_) );
  DFFR_X1 regBoiz_regfile_reg_4__16_ ( .D(n3998), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__16_) );
  DFFR_X1 regBoiz_regfile_reg_3__16_ ( .D(n3997), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__16_) );
  DFFR_X1 regBoiz_regfile_reg_2__16_ ( .D(n3996), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__16_) );
  DFFR_X1 regBoiz_regfile_reg_1__16_ ( .D(n3995), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__16_) );
  DFFR_X1 regBoiz_regfile_reg_0__16_ ( .D(n3994), .CK(clk), .RN(n6901), .Q(
        regBoiz_regfile_0__16_) );
  DFFR_X1 memBoi_memReg_22__regBoi_curData_reg ( .D(n3993), .CK(clk), .RN(
        n6874), .Q(wbBusWh[16]), .QN(n5654) );
  DFFR_X1 regBoiz_regfile_reg_31__15_ ( .D(n3992), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__15_) );
  DFFR_X1 regBoiz_regfile_reg_30__15_ ( .D(n3991), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__15_) );
  DFFR_X1 regBoiz_regfile_reg_29__15_ ( .D(n3990), .CK(clk), .RN(n6895), .Q(
        regBoiz_regfile_29__15_) );
  DFFR_X1 regBoiz_regfile_reg_28__15_ ( .D(n3989), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__15_) );
  DFFR_X1 regBoiz_regfile_reg_27__15_ ( .D(n3988), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_27__15_), .QN(n5544) );
  DFFR_X1 regBoiz_regfile_reg_25__15_ ( .D(n3986), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__15_), .QN(n5543) );
  DFFR_X1 regBoiz_regfile_reg_23__15_ ( .D(n3984), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__15_) );
  DFFR_X1 regBoiz_regfile_reg_22__15_ ( .D(n3983), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__15_) );
  DFFR_X1 regBoiz_regfile_reg_21__15_ ( .D(n3982), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_21__15_) );
  DFFR_X1 regBoiz_regfile_reg_20__15_ ( .D(n3981), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__15_) );
  DFFR_X1 regBoiz_regfile_reg_19__15_ ( .D(n3980), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_19__15_), .QN(n5542) );
  DFFR_X1 regBoiz_regfile_reg_17__15_ ( .D(n3978), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__15_), .QN(n5541) );
  DFFR_X1 regBoiz_regfile_reg_15__15_ ( .D(n3976), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__15_) );
  DFFR_X1 regBoiz_regfile_reg_14__15_ ( .D(n3975), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__15_) );
  DFFR_X1 regBoiz_regfile_reg_13__15_ ( .D(n3974), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_13__15_) );
  DFFR_X1 regBoiz_regfile_reg_12__15_ ( .D(n3973), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__15_) );
  DFFR_X1 regBoiz_regfile_reg_11__15_ ( .D(n3972), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__15_), .QN(n5540) );
  DFFR_X1 regBoiz_regfile_reg_10__15_ ( .D(n3971), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_10__15_), .QN(n5584) );
  DFFR_X1 regBoiz_regfile_reg_9__15_ ( .D(n3970), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_9__15_), .QN(n5539) );
  DFFR_X1 regBoiz_regfile_reg_8__15_ ( .D(n3969), .CK(clk), .RN(n6894), .Q(
        regBoiz_regfile_8__15_), .QN(n5420) );
  DFFR_X1 regBoiz_regfile_reg_7__15_ ( .D(n3968), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_7__15_) );
  DFFR_X1 regBoiz_regfile_reg_6__15_ ( .D(n3967), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_6__15_) );
  DFFR_X1 regBoiz_regfile_reg_5__15_ ( .D(n3966), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__15_) );
  DFFR_X1 regBoiz_regfile_reg_4__15_ ( .D(n3965), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__15_) );
  DFFR_X1 regBoiz_regfile_reg_3__15_ ( .D(n3964), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_3__15_), .QN(n5638) );
  DFFR_X1 regBoiz_regfile_reg_1__15_ ( .D(n3962), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__15_), .QN(n5538) );
  DFFR_X1 memBoi_memReg_23__regBoi_curData_reg ( .D(n3960), .CK(clk), .RN(
        n6900), .Q(wbBusWh[17]), .QN(n5653) );
  DFFR_X1 regBoiz_regfile_reg_31__14_ ( .D(n3959), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_31__14_) );
  DFFR_X1 regBoiz_regfile_reg_30__14_ ( .D(n3958), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__14_) );
  DFFR_X1 regBoiz_regfile_reg_29__14_ ( .D(n3957), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_29__14_) );
  DFFR_X1 regBoiz_regfile_reg_28__14_ ( .D(n3956), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__14_) );
  DFFR_X1 regBoiz_regfile_reg_27__14_ ( .D(n3955), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__14_), .QN(n5417) );
  DFFR_X1 regBoiz_regfile_reg_25__14_ ( .D(n3953), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__14_), .QN(n5416) );
  DFFR_X1 regBoiz_regfile_reg_24__14_ ( .D(n3952), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__14_), .QN(n5407) );
  DFFR_X1 regBoiz_regfile_reg_23__14_ ( .D(n3951), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_23__14_) );
  DFFR_X1 regBoiz_regfile_reg_22__14_ ( .D(n3950), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__14_) );
  DFFR_X1 regBoiz_regfile_reg_21__14_ ( .D(n3949), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__14_) );
  DFFR_X1 regBoiz_regfile_reg_20__14_ ( .D(n3948), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_20__14_) );
  DFFR_X1 regBoiz_regfile_reg_19__14_ ( .D(n3947), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__14_), .QN(n5415) );
  DFFR_X1 regBoiz_regfile_reg_17__14_ ( .D(n3945), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__14_), .QN(n5414) );
  DFFR_X1 regBoiz_regfile_reg_16__14_ ( .D(n3944), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__14_), .QN(n5406) );
  DFFR_X1 regBoiz_regfile_reg_15__14_ ( .D(n3943), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_15__14_) );
  DFFR_X1 regBoiz_regfile_reg_14__14_ ( .D(n3942), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__14_) );
  DFFR_X1 regBoiz_regfile_reg_13__14_ ( .D(n3941), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__14_) );
  DFFR_X1 regBoiz_regfile_reg_12__14_ ( .D(n3940), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_12__14_) );
  DFFR_X1 regBoiz_regfile_reg_11__14_ ( .D(n3939), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__14_), .QN(n5413) );
  DFFR_X1 regBoiz_regfile_reg_9__14_ ( .D(n3937), .CK(clk), .RN(n6896), .Q(
        regBoiz_regfile_9__14_), .QN(n5412) );
  DFFR_X1 regBoiz_regfile_reg_8__14_ ( .D(n3936), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_8__14_), .QN(n5405) );
  DFFR_X1 regBoiz_regfile_reg_7__14_ ( .D(n3935), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__14_) );
  DFFR_X1 regBoiz_regfile_reg_6__14_ ( .D(n3934), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__14_) );
  DFFR_X1 regBoiz_regfile_reg_5__14_ ( .D(n3933), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_5__14_) );
  DFFR_X1 regBoiz_regfile_reg_4__14_ ( .D(n3932), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__14_) );
  DFFR_X1 regBoiz_regfile_reg_3__14_ ( .D(n3931), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__14_), .QN(n5411) );
  DFFR_X1 regBoiz_regfile_reg_1__14_ ( .D(n3929), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__14_), .QN(n5410) );
  DFFR_X1 regBoiz_regfile_reg_0__14_ ( .D(n3928), .CK(clk), .RN(n6901), .Q(
        regBoiz_regfile_0__14_), .QN(n5404) );
  DFFR_X1 memBoi_memReg_24__regBoi_curData_reg ( .D(n3927), .CK(clk), .RN(
        n6874), .Q(wbBusWh[18]), .QN(n5652) );
  DFFR_X1 regBoiz_regfile_reg_29__13_ ( .D(n3924), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_29__13_) );
  DFFR_X1 regBoiz_regfile_reg_27__13_ ( .D(n3922), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_27__13_) );
  DFFR_X1 regBoiz_regfile_reg_26__13_ ( .D(n3921), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__13_) );
  DFFR_X1 regBoiz_regfile_reg_25__13_ ( .D(n3920), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__13_) );
  DFFR_X1 regBoiz_regfile_reg_24__13_ ( .D(n3919), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_24__13_) );
  DFFR_X1 regBoiz_regfile_reg_23__13_ ( .D(n3918), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__13_) );
  DFFR_X1 regBoiz_regfile_reg_22__13_ ( .D(n3917), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__13_) );
  DFFR_X1 regBoiz_regfile_reg_21__13_ ( .D(n3916), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_21__13_) );
  DFFR_X1 regBoiz_regfile_reg_20__13_ ( .D(n3915), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__13_) );
  DFFR_X1 regBoiz_regfile_reg_19__13_ ( .D(n3914), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_19__13_) );
  DFFR_X1 regBoiz_regfile_reg_18__13_ ( .D(n3913), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__13_) );
  DFFR_X1 regBoiz_regfile_reg_17__13_ ( .D(n3912), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__13_) );
  DFFR_X1 regBoiz_regfile_reg_16__13_ ( .D(n3911), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_16__13_) );
  DFFR_X1 regBoiz_regfile_reg_15__13_ ( .D(n3910), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__13_) );
  DFFR_X1 regBoiz_regfile_reg_14__13_ ( .D(n3909), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__13_) );
  DFFR_X1 regBoiz_regfile_reg_13__13_ ( .D(n3908), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_13__13_) );
  DFFR_X1 regBoiz_regfile_reg_12__13_ ( .D(n3907), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__13_) );
  DFFR_X1 regBoiz_regfile_reg_11__13_ ( .D(n3906), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__13_) );
  DFFR_X1 regBoiz_regfile_reg_10__13_ ( .D(n3905), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_10__13_) );
  DFFR_X1 regBoiz_regfile_reg_9__13_ ( .D(n3904), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_9__13_) );
  DFFR_X1 regBoiz_regfile_reg_8__13_ ( .D(n3903), .CK(clk), .RN(n6899), .Q(
        regBoiz_regfile_8__13_) );
  DFFR_X1 regBoiz_regfile_reg_7__13_ ( .D(n3902), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_7__13_) );
  DFFR_X1 regBoiz_regfile_reg_6__13_ ( .D(n3901), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_6__13_) );
  DFFR_X1 regBoiz_regfile_reg_5__13_ ( .D(n3900), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__13_) );
  DFFR_X1 regBoiz_regfile_reg_4__13_ ( .D(n3899), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__13_) );
  DFFR_X1 regBoiz_regfile_reg_3__13_ ( .D(n3898), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_3__13_) );
  DFFR_X1 regBoiz_regfile_reg_2__13_ ( .D(n3897), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_2__13_) );
  DFFR_X1 regBoiz_regfile_reg_1__13_ ( .D(n3896), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__13_) );
  DFFR_X1 regBoiz_regfile_reg_0__13_ ( .D(n3895), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__13_) );
  DFFR_X1 memBoi_memReg_25__regBoi_curData_reg ( .D(n3894), .CK(clk), .RN(
        n6900), .Q(wbBusWh[19]), .QN(n5651) );
  DFFR_X1 regBoiz_regfile_reg_31__12_ ( .D(n3893), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_31__12_) );
  DFFR_X1 regBoiz_regfile_reg_30__12_ ( .D(n3892), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__12_) );
  DFFR_X1 regBoiz_regfile_reg_29__12_ ( .D(n3891), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_29__12_) );
  DFFR_X1 regBoiz_regfile_reg_28__12_ ( .D(n3890), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__12_) );
  DFFR_X1 regBoiz_regfile_reg_27__12_ ( .D(n3889), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__12_) );
  DFFR_X1 regBoiz_regfile_reg_26__12_ ( .D(n3888), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_26__12_) );
  DFFR_X1 regBoiz_regfile_reg_25__12_ ( .D(n3887), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__12_) );
  DFFR_X1 regBoiz_regfile_reg_24__12_ ( .D(n3886), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__12_) );
  DFFR_X1 regBoiz_regfile_reg_23__12_ ( .D(n3885), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_23__12_) );
  DFFR_X1 regBoiz_regfile_reg_22__12_ ( .D(n3884), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__12_) );
  DFFR_X1 regBoiz_regfile_reg_21__12_ ( .D(n3883), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__12_) );
  DFFR_X1 regBoiz_regfile_reg_20__12_ ( .D(n3882), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_20__12_) );
  DFFR_X1 regBoiz_regfile_reg_19__12_ ( .D(n3881), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__12_) );
  DFFR_X1 regBoiz_regfile_reg_18__12_ ( .D(n3880), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_18__12_) );
  DFFR_X1 regBoiz_regfile_reg_17__12_ ( .D(n3879), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__12_) );
  DFFR_X1 regBoiz_regfile_reg_16__12_ ( .D(n3878), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__12_) );
  DFFR_X1 regBoiz_regfile_reg_13__12_ ( .D(n3875), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__12_) );
  DFFR_X1 regBoiz_regfile_reg_12__12_ ( .D(n3874), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_12__12_) );
  DFFR_X1 regBoiz_regfile_reg_11__12_ ( .D(n3873), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__12_) );
  DFFR_X1 regBoiz_regfile_reg_10__12_ ( .D(n3872), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__12_) );
  DFFR_X1 regBoiz_regfile_reg_9__12_ ( .D(n3871), .CK(clk), .RN(n6875), .Q(
        regBoiz_regfile_9__12_) );
  DFFR_X1 regBoiz_regfile_reg_8__12_ ( .D(n3870), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_8__12_) );
  DFFR_X1 regBoiz_regfile_reg_7__12_ ( .D(n3869), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__12_) );
  DFFR_X1 regBoiz_regfile_reg_6__12_ ( .D(n3868), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__12_) );
  DFFR_X1 regBoiz_regfile_reg_5__12_ ( .D(n3867), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_5__12_) );
  DFFR_X1 regBoiz_regfile_reg_4__12_ ( .D(n3866), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__12_) );
  DFFR_X1 regBoiz_regfile_reg_2__12_ ( .D(n3864), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__12_) );
  DFFR_X1 regBoiz_regfile_reg_0__12_ ( .D(n3862), .CK(clk), .RN(n6901), .Q(
        regBoiz_regfile_0__12_) );
  DFFR_X1 memBoi_memReg_26__regBoi_curData_reg ( .D(n3861), .CK(clk), .RN(
        n6874), .Q(wbBusWh[20]), .QN(n5650) );
  DFFR_X1 regBoiz_regfile_reg_31__11_ ( .D(n3860), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__11_) );
  DFFR_X1 regBoiz_regfile_reg_30__11_ ( .D(n3859), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__11_) );
  DFFR_X1 regBoiz_regfile_reg_29__11_ ( .D(n3858), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_29__11_) );
  DFFR_X1 regBoiz_regfile_reg_28__11_ ( .D(n3857), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__11_) );
  DFFR_X1 regBoiz_regfile_reg_27__11_ ( .D(n3856), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_27__11_) );
  DFFR_X1 regBoiz_regfile_reg_26__11_ ( .D(n3855), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__11_) );
  DFFR_X1 regBoiz_regfile_reg_25__11_ ( .D(n3854), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__11_) );
  DFFR_X1 regBoiz_regfile_reg_24__11_ ( .D(n3853), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_24__11_) );
  DFFR_X1 regBoiz_regfile_reg_23__11_ ( .D(n3852), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__11_) );
  DFFR_X1 regBoiz_regfile_reg_22__11_ ( .D(n3851), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__11_) );
  DFFR_X1 regBoiz_regfile_reg_21__11_ ( .D(n3850), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_21__11_) );
  DFFR_X1 regBoiz_regfile_reg_20__11_ ( .D(n3849), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__11_) );
  DFFR_X1 regBoiz_regfile_reg_19__11_ ( .D(n3848), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_19__11_) );
  DFFR_X1 regBoiz_regfile_reg_18__11_ ( .D(n3847), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__11_) );
  DFFR_X1 regBoiz_regfile_reg_17__11_ ( .D(n3846), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__11_) );
  DFFR_X1 regBoiz_regfile_reg_16__11_ ( .D(n3845), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_16__11_) );
  DFFR_X1 regBoiz_regfile_reg_15__11_ ( .D(n3844), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__11_) );
  DFFR_X1 regBoiz_regfile_reg_14__11_ ( .D(n3843), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__11_) );
  DFFR_X1 regBoiz_regfile_reg_13__11_ ( .D(n3842), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_13__11_) );
  DFFR_X1 regBoiz_regfile_reg_12__11_ ( .D(n3841), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__11_) );
  DFFR_X1 regBoiz_regfile_reg_11__11_ ( .D(n3840), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__11_) );
  DFFR_X1 regBoiz_regfile_reg_10__11_ ( .D(n3839), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_10__11_) );
  DFFR_X1 regBoiz_regfile_reg_9__11_ ( .D(n3838), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_9__11_) );
  DFFR_X1 regBoiz_regfile_reg_8__11_ ( .D(n3837), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_8__11_) );
  DFFR_X1 regBoiz_regfile_reg_7__11_ ( .D(n3836), .CK(clk), .RN(n6882), .Q(
        regBoiz_regfile_7__11_) );
  DFFR_X1 regBoiz_regfile_reg_6__11_ ( .D(n3835), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_6__11_) );
  DFFR_X1 regBoiz_regfile_reg_5__11_ ( .D(n3834), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__11_) );
  DFFR_X1 regBoiz_regfile_reg_4__11_ ( .D(n3833), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__11_) );
  DFFR_X1 regBoiz_regfile_reg_3__11_ ( .D(n3832), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_3__11_) );
  DFFR_X1 regBoiz_regfile_reg_2__11_ ( .D(n3831), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_2__11_) );
  DFFR_X1 regBoiz_regfile_reg_1__11_ ( .D(n3830), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__11_) );
  DFFR_X1 regBoiz_regfile_reg_0__11_ ( .D(n3829), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__11_) );
  DFFR_X1 memBoi_memReg_27__regBoi_curData_reg ( .D(n3828), .CK(clk), .RN(
        n6900), .Q(wbBusWh[21]), .QN(n5649) );
  DFFR_X1 regBoiz_regfile_reg_24__10_ ( .D(n3820), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__10_) );
  DFFR_X1 regBoiz_regfile_reg_20__10_ ( .D(n3816), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_20__10_) );
  DFFR_X1 regBoiz_regfile_reg_18__10_ ( .D(n3814), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_18__10_) );
  DFFR_X1 regBoiz_regfile_reg_17__10_ ( .D(n3813), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__10_) );
  DFFR_X1 regBoiz_regfile_reg_16__10_ ( .D(n3812), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__10_) );
  DFFR_X1 regBoiz_regfile_reg_13__10_ ( .D(n3809), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__10_) );
  DFFR_X1 regBoiz_regfile_reg_12__10_ ( .D(n3808), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_12__10_) );
  DFFR_X1 regBoiz_regfile_reg_10__10_ ( .D(n3806), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__10_) );
  DFFR_X1 regBoiz_regfile_reg_9__10_ ( .D(n3805), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_9__10_) );
  DFFR_X1 regBoiz_regfile_reg_8__10_ ( .D(n3804), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_8__10_) );
  DFFR_X1 regBoiz_regfile_reg_7__10_ ( .D(n3803), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__10_) );
  DFFR_X1 regBoiz_regfile_reg_6__10_ ( .D(n3802), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__10_) );
  DFFR_X1 regBoiz_regfile_reg_5__10_ ( .D(n3801), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_5__10_) );
  DFFR_X1 regBoiz_regfile_reg_4__10_ ( .D(n3800), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__10_) );
  DFFR_X1 regBoiz_regfile_reg_2__10_ ( .D(n3798), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__10_) );
  DFFR_X1 regBoiz_regfile_reg_1__10_ ( .D(n3797), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__10_) );
  DFFR_X1 regBoiz_regfile_reg_0__10_ ( .D(n3796), .CK(clk), .RN(n6901), .Q(
        regBoiz_regfile_0__10_) );
  DFFR_X1 memBoi_memReg_28__regBoi_curData_reg ( .D(n3795), .CK(clk), .RN(
        n6874), .Q(wbBusWh[22]), .QN(n5675) );
  DFFR_X1 regBoiz_regfile_reg_24__9_ ( .D(n3787), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_24__9_) );
  DFFR_X1 regBoiz_regfile_reg_18__9_ ( .D(n3781), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__9_) );
  DFFR_X1 regBoiz_regfile_reg_17__9_ ( .D(n3780), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__9_) );
  DFFR_X1 regBoiz_regfile_reg_16__9_ ( .D(n3779), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_16__9_) );
  DFFR_X1 regBoiz_regfile_reg_12__9_ ( .D(n3775), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__9_) );
  DFFR_X1 regBoiz_regfile_reg_11__9_ ( .D(n3774), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__9_) );
  DFFR_X1 regBoiz_regfile_reg_10__9_ ( .D(n3773), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_10__9_) );
  DFFR_X1 regBoiz_regfile_reg_8__9_ ( .D(n3771), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__9_) );
  DFFR_X1 regBoiz_regfile_reg_6__9_ ( .D(n3769), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_6__9_) );
  DFFR_X1 regBoiz_regfile_reg_5__9_ ( .D(n3768), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__9_) );
  DFFR_X1 regBoiz_regfile_reg_4__9_ ( .D(n3767), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__9_) );
  DFFR_X1 regBoiz_regfile_reg_3__9_ ( .D(n3766), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_3__9_) );
  DFFR_X1 regBoiz_regfile_reg_2__9_ ( .D(n3765), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_2__9_) );
  DFFR_X1 regBoiz_regfile_reg_1__9_ ( .D(n3764), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__9_) );
  DFFR_X1 regBoiz_regfile_reg_0__9_ ( .D(n3763), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__9_) );
  DFFR_X1 memBoi_memReg_29__regBoi_curData_reg ( .D(n3762), .CK(clk), .RN(
        n6900), .Q(wbBusWh[23]), .QN(n5674) );
  DFFR_X1 regBoiz_regfile_reg_30__8_ ( .D(n3760), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_30__8_) );
  DFFR_X1 regBoiz_regfile_reg_29__8_ ( .D(n3759), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__8_) );
  DFFR_X1 regBoiz_regfile_reg_28__8_ ( .D(n3758), .CK(clk), .RN(n6889), .Q(
        regBoiz_regfile_28__8_) );
  DFFR_X1 regBoiz_regfile_reg_27__8_ ( .D(n3757), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__8_) );
  DFFR_X1 regBoiz_regfile_reg_26__8_ ( .D(n3756), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__8_) );
  DFFR_X1 regBoiz_regfile_reg_25__8_ ( .D(n3755), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_25__8_) );
  DFFR_X1 regBoiz_regfile_reg_24__8_ ( .D(n3754), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__8_) );
  DFFR_X1 regBoiz_regfile_reg_22__8_ ( .D(n3752), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_22__8_) );
  DFFR_X1 regBoiz_regfile_reg_21__8_ ( .D(n3751), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__8_) );
  DFFR_X1 regBoiz_regfile_reg_20__8_ ( .D(n3750), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__8_) );
  DFFR_X1 regBoiz_regfile_reg_19__8_ ( .D(n3749), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__8_) );
  DFFR_X1 regBoiz_regfile_reg_18__8_ ( .D(n3748), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__8_) );
  DFFR_X1 regBoiz_regfile_reg_17__8_ ( .D(n3747), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_17__8_) );
  DFFR_X1 regBoiz_regfile_reg_16__8_ ( .D(n3746), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__8_) );
  DFFR_X1 regBoiz_regfile_reg_14__8_ ( .D(n3744), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_14__8_) );
  DFFR_X1 regBoiz_regfile_reg_13__8_ ( .D(n3743), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__8_) );
  DFFR_X1 regBoiz_regfile_reg_12__8_ ( .D(n3742), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__8_) );
  DFFR_X1 regBoiz_regfile_reg_11__8_ ( .D(n3741), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_11__8_) );
  DFFR_X1 regBoiz_regfile_reg_10__8_ ( .D(n3740), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__8_) );
  DFFR_X1 regBoiz_regfile_reg_9__8_ ( .D(n3739), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_9__8_) );
  DFFR_X1 regBoiz_regfile_reg_8__8_ ( .D(n3738), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_8__8_) );
  DFFR_X1 regBoiz_regfile_reg_7__8_ ( .D(n3737), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_7__8_) );
  DFFR_X1 regBoiz_regfile_reg_6__8_ ( .D(n3736), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__8_) );
  DFFR_X1 regBoiz_regfile_reg_5__8_ ( .D(n3735), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__8_) );
  DFFR_X1 regBoiz_regfile_reg_4__8_ ( .D(n3734), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_4__8_) );
  DFFR_X1 regBoiz_regfile_reg_3__8_ ( .D(n3733), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__8_) );
  DFFR_X1 regBoiz_regfile_reg_2__8_ ( .D(n3732), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__8_) );
  DFFR_X1 regBoiz_regfile_reg_1__8_ ( .D(n3731), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_1__8_) );
  DFFR_X1 regBoiz_regfile_reg_0__8_ ( .D(n3730), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__8_) );
  DFFR_X1 memBoi_memReg_30__regBoi_curData_reg ( .D(n3729), .CK(clk), .RN(
        n6901), .Q(wbBusWh[24]), .QN(n5673) );
  DFFR_X1 regBoiz_regfile_reg_31__7_ ( .D(n3728), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__7_) );
  DFFR_X1 regBoiz_regfile_reg_30__7_ ( .D(n3727), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__7_) );
  DFFR_X1 regBoiz_regfile_reg_29__7_ ( .D(n3726), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__7_) );
  DFFR_X1 regBoiz_regfile_reg_28__7_ ( .D(n3725), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__7_) );
  DFFR_X1 regBoiz_regfile_reg_27__7_ ( .D(n3724), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_27__7_) );
  DFFR_X1 regBoiz_regfile_reg_26__7_ ( .D(n3723), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__7_) );
  DFFR_X1 regBoiz_regfile_reg_25__7_ ( .D(n3722), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__7_) );
  DFFR_X1 regBoiz_regfile_reg_24__7_ ( .D(n3721), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_24__7_) );
  DFFR_X1 regBoiz_regfile_reg_23__7_ ( .D(n3720), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__7_) );
  DFFR_X1 regBoiz_regfile_reg_22__7_ ( .D(n3719), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__7_) );
  DFFR_X1 regBoiz_regfile_reg_21__7_ ( .D(n3718), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_21__7_) );
  DFFR_X1 regBoiz_regfile_reg_20__7_ ( .D(n3717), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__7_) );
  DFFR_X1 regBoiz_regfile_reg_19__7_ ( .D(n3716), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_19__7_) );
  DFFR_X1 regBoiz_regfile_reg_18__7_ ( .D(n3715), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__7_) );
  DFFR_X1 regBoiz_regfile_reg_17__7_ ( .D(n3714), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__7_) );
  DFFR_X1 regBoiz_regfile_reg_16__7_ ( .D(n3713), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_16__7_) );
  DFFR_X1 regBoiz_regfile_reg_12__7_ ( .D(n3709), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__7_) );
  DFFR_X1 regBoiz_regfile_reg_10__7_ ( .D(n3707), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_10__7_) );
  DFFR_X1 regBoiz_regfile_reg_9__7_ ( .D(n3706), .CK(clk), .RN(n6943), .Q(
        regBoiz_regfile_9__7_) );
  DFFR_X1 regBoiz_regfile_reg_8__7_ ( .D(n3705), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__7_) );
  DFFR_X1 regBoiz_regfile_reg_6__7_ ( .D(n3703), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_6__7_) );
  DFFR_X1 regBoiz_regfile_reg_5__7_ ( .D(n3702), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__7_) );
  DFFR_X1 regBoiz_regfile_reg_4__7_ ( .D(n3701), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__7_) );
  DFFR_X1 regBoiz_regfile_reg_3__7_ ( .D(n3700), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_3__7_) );
  DFFR_X1 regBoiz_regfile_reg_2__7_ ( .D(n3699), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_2__7_) );
  DFFR_X1 regBoiz_regfile_reg_1__7_ ( .D(n3698), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__7_) );
  DFFR_X1 regBoiz_regfile_reg_0__7_ ( .D(n3697), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__7_) );
  DFFR_X1 memBoi_memReg_31__regBoi_curData_reg ( .D(n3696), .CK(clk), .RN(
        n6874), .Q(wbBusWh[25]), .QN(n5684) );
  DFFR_X1 regBoiz_regfile_reg_30__6_ ( .D(n3694), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_30__6_) );
  DFFR_X1 regBoiz_regfile_reg_29__6_ ( .D(n3693), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__6_) );
  DFFR_X1 regBoiz_regfile_reg_28__6_ ( .D(n3692), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_28__6_) );
  DFFR_X1 regBoiz_regfile_reg_27__6_ ( .D(n3691), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__6_) );
  DFFR_X1 regBoiz_regfile_reg_26__6_ ( .D(n3690), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__6_) );
  DFFR_X1 regBoiz_regfile_reg_25__6_ ( .D(n3689), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_25__6_) );
  DFFR_X1 regBoiz_regfile_reg_24__6_ ( .D(n3688), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__6_) );
  DFFR_X1 regBoiz_regfile_reg_23__6_ ( .D(n3687), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__6_) );
  DFFR_X1 regBoiz_regfile_reg_22__6_ ( .D(n3686), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_22__6_) );
  DFFR_X1 regBoiz_regfile_reg_21__6_ ( .D(n3685), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__6_) );
  DFFR_X1 regBoiz_regfile_reg_20__6_ ( .D(n3684), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__6_) );
  DFFR_X1 regBoiz_regfile_reg_19__6_ ( .D(n3683), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__6_) );
  DFFR_X1 regBoiz_regfile_reg_18__6_ ( .D(n3682), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__6_) );
  DFFR_X1 regBoiz_regfile_reg_17__6_ ( .D(n3681), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_17__6_) );
  DFFR_X1 regBoiz_regfile_reg_16__6_ ( .D(n3680), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__6_) );
  DFFR_X1 regBoiz_regfile_reg_14__6_ ( .D(n3678), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_14__6_) );
  DFFR_X1 regBoiz_regfile_reg_13__6_ ( .D(n3677), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__6_) );
  DFFR_X1 regBoiz_regfile_reg_12__6_ ( .D(n3676), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__6_) );
  DFFR_X1 regBoiz_regfile_reg_11__6_ ( .D(n3675), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_11__6_) );
  DFFR_X1 regBoiz_regfile_reg_10__6_ ( .D(n3674), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__6_) );
  DFFR_X1 regBoiz_regfile_reg_9__6_ ( .D(n3673), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_9__6_) );
  DFFR_X1 regBoiz_regfile_reg_8__6_ ( .D(n3672), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_8__6_) );
  DFFR_X1 regBoiz_regfile_reg_7__6_ ( .D(n3671), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_7__6_) );
  DFFR_X1 regBoiz_regfile_reg_6__6_ ( .D(n3670), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__6_) );
  DFFR_X1 regBoiz_regfile_reg_5__6_ ( .D(n3669), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__6_) );
  DFFR_X1 regBoiz_regfile_reg_4__6_ ( .D(n3668), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_4__6_) );
  DFFR_X1 regBoiz_regfile_reg_3__6_ ( .D(n3667), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__6_) );
  DFFR_X1 regBoiz_regfile_reg_2__6_ ( .D(n3666), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__6_) );
  DFFR_X1 regBoiz_regfile_reg_1__6_ ( .D(n3665), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_1__6_) );
  DFFR_X1 regBoiz_regfile_reg_0__6_ ( .D(n3664), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__6_) );
  DFFR_X1 memBoi_memReg_32__regBoi_curData_reg ( .D(n3663), .CK(clk), .RN(
        n6901), .Q(wbBusWh[26]), .QN(n5672) );
  DFFR_X1 regBoiz_regfile_reg_31__5_ ( .D(n3662), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__5_) );
  DFFR_X1 regBoiz_regfile_reg_30__5_ ( .D(n3661), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__5_) );
  DFFR_X1 regBoiz_regfile_reg_28__5_ ( .D(n3659), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__5_) );
  DFFR_X1 regBoiz_regfile_reg_27__5_ ( .D(n3658), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_27__5_) );
  DFFR_X1 regBoiz_regfile_reg_26__5_ ( .D(n3657), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__5_) );
  DFFR_X1 regBoiz_regfile_reg_25__5_ ( .D(n3656), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__5_) );
  DFFR_X1 regBoiz_regfile_reg_24__5_ ( .D(n3655), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_24__5_) );
  DFFR_X1 regBoiz_regfile_reg_23__5_ ( .D(n3654), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__5_) );
  DFFR_X1 regBoiz_regfile_reg_22__5_ ( .D(n3653), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__5_) );
  DFFR_X1 regBoiz_regfile_reg_21__5_ ( .D(n3652), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_21__5_) );
  DFFR_X1 regBoiz_regfile_reg_20__5_ ( .D(n3651), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__5_) );
  DFFR_X1 regBoiz_regfile_reg_19__5_ ( .D(n3650), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_19__5_) );
  DFFR_X1 regBoiz_regfile_reg_18__5_ ( .D(n3649), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__5_) );
  DFFR_X1 regBoiz_regfile_reg_17__5_ ( .D(n3648), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__5_) );
  DFFR_X1 regBoiz_regfile_reg_16__5_ ( .D(n3647), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_16__5_) );
  DFFR_X1 regBoiz_regfile_reg_15__5_ ( .D(n3646), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__5_) );
  DFFR_X1 regBoiz_regfile_reg_14__5_ ( .D(n3645), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__5_) );
  DFFR_X1 regBoiz_regfile_reg_13__5_ ( .D(n3644), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_13__5_) );
  DFFR_X1 regBoiz_regfile_reg_12__5_ ( .D(n3643), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__5_) );
  DFFR_X1 regBoiz_regfile_reg_11__5_ ( .D(n3642), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__5_) );
  DFFR_X1 regBoiz_regfile_reg_10__5_ ( .D(n3641), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_10__5_) );
  DFFR_X1 regBoiz_regfile_reg_9__5_ ( .D(n3640), .CK(clk), .RN(n6943), .Q(
        regBoiz_regfile_9__5_) );
  DFFR_X1 regBoiz_regfile_reg_8__5_ ( .D(n3639), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__5_) );
  DFFR_X1 regBoiz_regfile_reg_7__5_ ( .D(n3638), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__5_) );
  DFFR_X1 regBoiz_regfile_reg_6__5_ ( .D(n3637), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_6__5_) );
  DFFR_X1 regBoiz_regfile_reg_5__5_ ( .D(n3636), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__5_) );
  DFFR_X1 regBoiz_regfile_reg_4__5_ ( .D(n3635), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__5_) );
  DFFR_X1 regBoiz_regfile_reg_3__5_ ( .D(n3634), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_3__5_) );
  DFFR_X1 regBoiz_regfile_reg_2__5_ ( .D(n3633), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_2__5_) );
  DFFR_X1 regBoiz_regfile_reg_1__5_ ( .D(n3632), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__5_) );
  DFFR_X1 regBoiz_regfile_reg_0__5_ ( .D(n3631), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__5_) );
  DFFR_X1 memBoi_memReg_33__regBoi_curData_reg ( .D(n3630), .CK(clk), .RN(
        n6874), .Q(wbBusWh[27]), .QN(n5688) );
  DFFR_X1 regBoiz_regfile_reg_24__4_ ( .D(n3622), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__4_) );
  DFFR_X1 regBoiz_regfile_reg_18__4_ ( .D(n3616), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__4_), .QN(n6352) );
  DFFR_X1 regBoiz_regfile_reg_16__4_ ( .D(n3614), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__4_) );
  DFFR_X1 regBoiz_regfile_reg_8__4_ ( .D(n3606), .CK(clk), .RN(n6883), .Q(
        regBoiz_regfile_8__4_), .QN(n6253) );
  DFFR_X1 regBoiz_regfile_reg_4__4_ ( .D(n3602), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_4__4_) );
  DFFR_X1 regBoiz_regfile_reg_2__4_ ( .D(n3600), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__4_) );
  DFFR_X1 regBoiz_regfile_reg_1__4_ ( .D(n3599), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_1__4_) );
  DFFR_X1 regBoiz_regfile_reg_0__4_ ( .D(n3598), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__4_), .QN(n6254) );
  DFFR_X1 memBoi_memReg_34__regBoi_curData_reg ( .D(n3597), .CK(clk), .RN(
        n6901), .Q(wbBusWh[28]), .QN(n5671) );
  DFFR_X1 regBoiz_regfile_reg_28__3_ ( .D(n3593), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__3_) );
  DFFR_X1 regBoiz_regfile_reg_26__3_ ( .D(n3591), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__3_) );
  DFFR_X1 regBoiz_regfile_reg_25__3_ ( .D(n3590), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__3_) );
  DFFR_X1 regBoiz_regfile_reg_24__3_ ( .D(n3589), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_24__3_) );
  DFFR_X1 regBoiz_regfile_reg_22__3_ ( .D(n3587), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__3_) );
  DFFR_X1 regBoiz_regfile_reg_21__3_ ( .D(n3586), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_21__3_), .QN(n6256) );
  DFFR_X1 regBoiz_regfile_reg_20__3_ ( .D(n3585), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__3_) );
  DFFR_X1 regBoiz_regfile_reg_19__3_ ( .D(n3584), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_19__3_) );
  DFFR_X1 regBoiz_regfile_reg_18__3_ ( .D(n3583), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__3_) );
  DFFR_X1 regBoiz_regfile_reg_17__3_ ( .D(n3582), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_17__3_) );
  DFFR_X1 regBoiz_regfile_reg_16__3_ ( .D(n3581), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_16__3_) );
  DFFR_X1 regBoiz_regfile_reg_13__3_ ( .D(n3578), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_13__3_) );
  DFFR_X1 regBoiz_regfile_reg_12__3_ ( .D(n3577), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__3_) );
  DFFR_X1 regBoiz_regfile_reg_11__3_ ( .D(n3576), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__3_) );
  DFFR_X1 regBoiz_regfile_reg_10__3_ ( .D(n3575), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_10__3_) );
  DFFR_X1 regBoiz_regfile_reg_9__3_ ( .D(n3574), .CK(clk), .RN(n6943), .Q(
        regBoiz_regfile_9__3_) );
  DFFR_X1 regBoiz_regfile_reg_8__3_ ( .D(n3573), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__3_) );
  DFFR_X1 regBoiz_regfile_reg_7__3_ ( .D(n3572), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__3_) );
  DFFR_X1 regBoiz_regfile_reg_6__3_ ( .D(n3571), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_6__3_) );
  DFFR_X1 regBoiz_regfile_reg_5__3_ ( .D(n3570), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__3_) );
  DFFR_X1 regBoiz_regfile_reg_4__3_ ( .D(n3569), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_4__3_) );
  DFFR_X1 regBoiz_regfile_reg_3__3_ ( .D(n3568), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_3__3_) );
  DFFR_X1 regBoiz_regfile_reg_2__3_ ( .D(n3567), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_2__3_) );
  DFFR_X1 regBoiz_regfile_reg_1__3_ ( .D(n3566), .CK(clk), .RN(n6917), .Q(
        regBoiz_regfile_1__3_) );
  DFFR_X1 regBoiz_regfile_reg_0__3_ ( .D(n3565), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__3_) );
  DFFR_X1 memBoi_memReg_35__regBoi_curData_reg ( .D(n3564), .CK(clk), .RN(
        n6874), .Q(wbBusWh[29]), .QN(n5669) );
  DFFR_X1 regBoiz_regfile_reg_30__2_ ( .D(n3562), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__2_) );
  DFFR_X1 regBoiz_regfile_reg_29__2_ ( .D(n3561), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__2_) );
  DFFR_X1 regBoiz_regfile_reg_28__2_ ( .D(n3560), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__2_) );
  DFFR_X1 regBoiz_regfile_reg_27__2_ ( .D(n3559), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__2_) );
  DFFR_X1 regBoiz_regfile_reg_26__2_ ( .D(n3558), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__2_) );
  DFFR_X1 regBoiz_regfile_reg_25__2_ ( .D(n3557), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__2_) );
  DFFR_X1 regBoiz_regfile_reg_24__2_ ( .D(n3556), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__2_) );
  DFFR_X1 regBoiz_regfile_reg_23__2_ ( .D(n3555), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__2_) );
  DFFR_X1 regBoiz_regfile_reg_22__2_ ( .D(n3554), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__2_) );
  DFFR_X1 regBoiz_regfile_reg_21__2_ ( .D(n3553), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__2_) );
  DFFR_X1 regBoiz_regfile_reg_20__2_ ( .D(n3552), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__2_) );
  DFFR_X1 regBoiz_regfile_reg_19__2_ ( .D(n3551), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__2_) );
  DFFR_X1 regBoiz_regfile_reg_18__2_ ( .D(n3550), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__2_) );
  DFFR_X1 regBoiz_regfile_reg_17__2_ ( .D(n3549), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__2_) );
  DFFR_X1 regBoiz_regfile_reg_16__2_ ( .D(n3548), .CK(clk), .RN(n6863), .Q(
        regBoiz_regfile_16__2_) );
  DFFR_X1 regBoiz_regfile_reg_15__2_ ( .D(n3547), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__2_) );
  DFFR_X1 regBoiz_regfile_reg_14__2_ ( .D(n3546), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__2_) );
  DFFR_X1 regBoiz_regfile_reg_13__2_ ( .D(n3545), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__2_) );
  DFFR_X1 regBoiz_regfile_reg_12__2_ ( .D(n3544), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__2_) );
  DFFR_X1 regBoiz_regfile_reg_11__2_ ( .D(n3543), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__2_) );
  DFFR_X1 regBoiz_regfile_reg_10__2_ ( .D(n3542), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__2_) );
  DFFR_X1 regBoiz_regfile_reg_9__2_ ( .D(n3541), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_9__2_) );
  DFFR_X1 regBoiz_regfile_reg_8__2_ ( .D(n3540), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_8__2_) );
  DFFR_X1 regBoiz_regfile_reg_7__2_ ( .D(n3539), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_7__2_) );
  DFFR_X1 regBoiz_regfile_reg_6__2_ ( .D(n3538), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__2_) );
  DFFR_X1 regBoiz_regfile_reg_5__2_ ( .D(n3537), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__2_) );
  DFFR_X1 regBoiz_regfile_reg_4__2_ ( .D(n3536), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__2_) );
  DFFR_X1 regBoiz_regfile_reg_3__2_ ( .D(n3535), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__2_) );
  DFFR_X1 regBoiz_regfile_reg_2__2_ ( .D(n3534), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__2_) );
  DFFR_X1 regBoiz_regfile_reg_1__2_ ( .D(n3533), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__2_) );
  DFFR_X1 regBoiz_regfile_reg_0__2_ ( .D(n3532), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_0__2_) );
  DFFR_X1 memBoi_memReg_36__regBoi_curData_reg ( .D(n3531), .CK(clk), .RN(
        n6901), .Q(wbBusWh[30]), .QN(n5659) );
  DFFR_X1 regBoiz_regfile_reg_27__1_ ( .D(n3526), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__1_) );
  DFFR_X1 regBoiz_regfile_reg_26__1_ ( .D(n3525), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__1_) );
  DFFR_X1 regBoiz_regfile_reg_25__1_ ( .D(n3524), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__1_) );
  DFFR_X1 regBoiz_regfile_reg_24__1_ ( .D(n3523), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__1_) );
  DFFR_X1 regBoiz_regfile_reg_23__1_ ( .D(n3522), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__1_) );
  DFFR_X1 regBoiz_regfile_reg_22__1_ ( .D(n3521), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__1_) );
  DFFR_X1 regBoiz_regfile_reg_21__1_ ( .D(n3520), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__1_) );
  DFFR_X1 regBoiz_regfile_reg_20__1_ ( .D(n3519), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__1_) );
  DFFR_X1 regBoiz_regfile_reg_19__1_ ( .D(n3518), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__1_) );
  DFFR_X1 regBoiz_regfile_reg_18__1_ ( .D(n3517), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__1_) );
  DFFR_X1 regBoiz_regfile_reg_17__1_ ( .D(n3516), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__1_) );
  DFFR_X1 regBoiz_regfile_reg_16__1_ ( .D(n3515), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__1_) );
  DFFR_X1 regBoiz_regfile_reg_15__1_ ( .D(n3514), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__1_) );
  DFFR_X1 regBoiz_regfile_reg_14__1_ ( .D(n3513), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__1_) );
  DFFR_X1 regBoiz_regfile_reg_13__1_ ( .D(n3512), .CK(clk), .RN(n6907), .Q(
        regBoiz_regfile_13__1_) );
  DFFR_X1 regBoiz_regfile_reg_12__1_ ( .D(n3511), .CK(clk), .RN(n6906), .Q(
        regBoiz_regfile_12__1_) );
  DFFR_X1 regBoiz_regfile_reg_11__1_ ( .D(n3510), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__1_) );
  DFFR_X1 regBoiz_regfile_reg_10__1_ ( .D(n3509), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__1_) );
  DFFR_X1 regBoiz_regfile_reg_9__1_ ( .D(n3508), .CK(clk), .RN(n6874), .Q(
        regBoiz_regfile_9__1_) );
  DFFR_X1 regBoiz_regfile_reg_8__1_ ( .D(n3507), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__1_) );
  DFFR_X1 regBoiz_regfile_reg_6__1_ ( .D(n3505), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__1_) );
  DFFR_X1 regBoiz_regfile_reg_5__1_ ( .D(n3504), .CK(clk), .RN(n6938), .Q(
        regBoiz_regfile_5__1_) );
  DFFR_X1 regBoiz_regfile_reg_4__1_ ( .D(n3503), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_4__1_) );
  DFFR_X1 regBoiz_regfile_reg_3__1_ ( .D(n3502), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__1_) );
  DFFR_X1 regBoiz_regfile_reg_2__1_ ( .D(n3501), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__1_) );
  DFFR_X1 regBoiz_regfile_reg_1__1_ ( .D(n3500), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__1_) );
  DFFR_X1 regBoiz_regfile_reg_0__1_ ( .D(n3499), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__1_) );
  DFFR_X1 memBoi_memReg_37__regBoi_curData_reg ( .D(n3498), .CK(clk), .RN(
        n6873), .Q(wbBusWh[31]), .QN(n5648) );
  DFFR_X1 regBoiz_regfile_reg_31__0_ ( .D(n3497), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__0_) );
  DFFR_X1 regBoiz_regfile_reg_30__0_ ( .D(n3496), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__0_) );
  DFFR_X1 regBoiz_regfile_reg_29__0_ ( .D(n3495), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_29__0_) );
  DFFR_X1 regBoiz_regfile_reg_28__0_ ( .D(n3494), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__0_) );
  DFFR_X1 regBoiz_regfile_reg_27__0_ ( .D(n3493), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_27__0_) );
  DFFR_X1 regBoiz_regfile_reg_26__0_ ( .D(n3492), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__0_) );
  DFFR_X1 regBoiz_regfile_reg_25__0_ ( .D(n3491), .CK(clk), .RN(n6850), .Q(
        regBoiz_regfile_25__0_) );
  DFFR_X1 regBoiz_regfile_reg_24__0_ ( .D(n3490), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_24__0_) );
  DFFR_X1 regBoiz_regfile_reg_23__0_ ( .D(n3489), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_23__0_) );
  DFFR_X1 regBoiz_regfile_reg_22__0_ ( .D(n3488), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__0_) );
  DFFR_X1 regBoiz_regfile_reg_21__0_ ( .D(n3487), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_21__0_) );
  DFFR_X1 regBoiz_regfile_reg_20__0_ ( .D(n3486), .CK(clk), .RN(n6857), .Q(
        regBoiz_regfile_20__0_) );
  DFFR_X1 regBoiz_regfile_reg_19__0_ ( .D(n3485), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_19__0_) );
  DFFR_X1 regBoiz_regfile_reg_18__0_ ( .D(n3484), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__0_) );
  DFFR_X1 regBoiz_regfile_reg_17__0_ ( .D(n3483), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__0_) );
  DFFR_X1 regBoiz_regfile_reg_16__0_ ( .D(n3482), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_16__0_) );
  DFFR_X1 regBoiz_regfile_reg_15__0_ ( .D(n3481), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__0_) );
  DFFR_X1 regBoiz_regfile_reg_14__0_ ( .D(n3480), .CK(clk), .RN(n6866), .Q(
        regBoiz_regfile_14__0_) );
  DFFR_X1 regBoiz_regfile_reg_13__0_ ( .D(n3479), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_13__0_) );
  DFFR_X1 regBoiz_regfile_reg_12__0_ ( .D(n3478), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_12__0_) );
  DFFR_X1 regBoiz_regfile_reg_11__0_ ( .D(n3477), .CK(clk), .RN(n6870), .Q(
        regBoiz_regfile_11__0_) );
  DFFR_X1 regBoiz_regfile_reg_10__0_ ( .D(n3476), .CK(clk), .RN(n6872), .Q(
        regBoiz_regfile_10__0_) );
  DFFR_X1 regBoiz_regfile_reg_9__0_ ( .D(n3475), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_9__0_) );
  DFFR_X1 regBoiz_regfile_reg_8__0_ ( .D(n3474), .CK(clk), .RN(n6877), .Q(
        regBoiz_regfile_8__0_) );
  DFFR_X1 regBoiz_regfile_reg_7__0_ ( .D(n3473), .CK(clk), .RN(n6936), .Q(
        regBoiz_regfile_7__0_) );
  DFFR_X1 regBoiz_regfile_reg_6__0_ ( .D(n3472), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_6__0_) );
  DFFR_X1 regBoiz_regfile_reg_5__0_ ( .D(n3471), .CK(clk), .RN(n6838), .Q(
        regBoiz_regfile_5__0_) );
  DFFR_X1 regBoiz_regfile_reg_4__0_ ( .D(n3470), .CK(clk), .RN(n6839), .Q(
        regBoiz_regfile_4__0_) );
  DFFR_X1 regBoiz_regfile_reg_3__0_ ( .D(n3469), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_3__0_) );
  DFFR_X1 regBoiz_regfile_reg_2__0_ ( .D(n3468), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_2__0_) );
  DFFR_X1 regBoiz_regfile_reg_1__0_ ( .D(n3467), .CK(clk), .RN(n6858), .Q(
        regBoiz_regfile_1__0_) );
  DFFR_X1 regBoiz_regfile_reg_0__0_ ( .D(n3466), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__0_) );
  DFF_X2 aluBoi_multBoi_count_reg_0_ ( .D(aluBoi_multBoi_N71), .CK(clk), .Q(
        aluBoi_multBoi_count_0_) );
  DFF_X2 aluBoi_multBoi_count_reg_1_ ( .D(aluBoi_multBoi_N72), .CK(clk), .Q(
        aluBoi_multBoi_count_1_) );
  DFF_X2 aluBoi_multBoi_count_reg_2_ ( .D(aluBoi_multBoi_N73), .CK(clk), .Q(
        aluBoi_multBoi_count_2_) );
  DFF_X2 aluBoi_multBoi_runProd_reg_64_ ( .D(aluBoi_multBoi_N70), .CK(clk), 
        .Q(net129670) );
  DFF_X2 aluBoi_multBoi_runProd_reg_58_ ( .D(aluBoi_multBoi_N64), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[54]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_38_ ( .D(aluBoi_multBoi_N44), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[34]), .QN(n5552) );
  DFF_X2 aluBoi_multBoi_runProd_reg_34_ ( .D(aluBoi_multBoi_N40), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[30]), .QN(n5678) );
  DFF_X2 aluBoi_multBoi_runProd_reg_30_ ( .D(aluBoi_multBoi_N36), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[26]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_35_ ( .D(aluBoi_multBoi_N41), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[31]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_31_ ( .D(aluBoi_multBoi_N37), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[27]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_27_ ( .D(n13679), .CK(clk), .Q(
        aluBoi_multBoi_temppp[23]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_53_ ( .D(aluBoi_multBoi_N59), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[49]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_33_ ( .D(n5036), .CK(clk), .Q(
        aluBoi_multBoi_temppp[29]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_29_ ( .D(aluBoi_multBoi_N35), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[25]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_25_ ( .D(n13681), .CK(clk), .Q(
        aluBoi_multBoi_temppp[21]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_26_ ( .D(n13678), .CK(clk), .Q(
        aluBoi_multBoi_temppp[22]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_52_ ( .D(aluBoi_multBoi_N58), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[48]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_48_ ( .D(aluBoi_multBoi_N54), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[44]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_36_ ( .D(aluBoi_multBoi_N42), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[32]), .QN(n5679) );
  DFF_X2 aluBoi_multBoi_runProd_reg_32_ ( .D(aluBoi_multBoi_N38), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[28]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_28_ ( .D(aluBoi_multBoi_N34), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[24]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_24_ ( .D(n13684), .CK(clk), .Q(
        aluBoi_multBoi_temppp[20]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_23_ ( .D(n13680), .CK(clk), .Q(
        aluBoi_multBoi_temppp[19]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_22_ ( .D(n13683), .CK(clk), .Q(
        aluBoi_multBoi_temppp[18]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_21_ ( .D(n13682), .CK(clk), .Q(
        aluBoi_multBoi_temppp[17]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_17_ ( .D(n13688), .CK(clk), .Q(
        aluBoi_multBoi_temppp[13]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_18_ ( .D(n13687), .CK(clk), .Q(
        aluBoi_multBoi_temppp[14]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_19_ ( .D(n13686), .CK(clk), .Q(
        aluBoi_multBoi_temppp[15]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_20_ ( .D(n13685), .CK(clk), .Q(
        aluBoi_multBoi_temppp[16]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_16_ ( .D(n13692), .CK(clk), .Q(
        aluBoi_multBoi_temppp[12]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_12_ ( .D(n13693), .CK(clk), .Q(
        aluBoi_multBoi_temppp[8]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_13_ ( .D(n13689), .CK(clk), .Q(
        aluBoi_multBoi_temppp[9]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_14_ ( .D(n13690), .CK(clk), .Q(
        aluBoi_multBoi_temppp[10]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_15_ ( .D(n13691), .CK(clk), .Q(
        aluBoi_multBoi_temppp[11]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_11_ ( .D(n13697), .CK(clk), .Q(
        aluBoi_multBoi_temppp[7]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_7_ ( .D(n13698), .CK(clk), .Q(
        aluBoi_multBoi_temppp[3]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_3_ ( .D(n13699), .CK(clk), .Q(
        aluBoi_multOut[2]), .QN(n5304) );
  DFF_X2 aluBoi_multBoi_runProd_reg_8_ ( .D(n13694), .CK(clk), .Q(
        aluBoi_multBoi_temppp[4]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_4_ ( .D(n13700), .CK(clk), .Q(
        aluBoi_multBoi_temppp[0]), .QN(n5471) );
  DFF_X2 aluBoi_multBoi_runProd_reg_0_ ( .D(aluBoi_multBoi_N6), .CK(clk), .Q(
        aluBoi_multBoi_runProd_0_), .QN(n5690) );
  DFF_X2 aluBoi_multBoi_runProd_reg_9_ ( .D(n13695), .CK(clk), .Q(
        aluBoi_multBoi_temppp[5]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_5_ ( .D(n13701), .CK(clk), .Q(
        aluBoi_multBoi_temppp[1]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_1_ ( .D(n13702), .CK(clk), .Q(
        aluBoi_multOut[0]), .QN(n5307) );
  DFF_X2 aluBoi_multBoi_runProd_reg_10_ ( .D(n13696), .CK(clk), .Q(
        aluBoi_multBoi_temppp[6]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_6_ ( .D(n13703), .CK(clk), .Q(
        aluBoi_multBoi_temppp[2]) );
  DFF_X2 aluBoi_multBoi_runProd_reg_2_ ( .D(n13704), .CK(clk), .Q(
        aluBoi_multOut[1]), .QN(n5319) );
  DLH_X2 aluBoi_condBoi_outBit_reg ( .G(aluBoi_condBoi_N24), .D(
        aluBoi_condBoi_N25), .Q(aluBoi_condOut_0_) );
  DFF_X2 aluBoi_multBoi_ready_reg ( .D(n4873), .CK(clk), .QN(n5691) );
  DFFRS_X2 ifBoi_pcOut_reg_0_ ( .D(n4713), .CK(clk), .RN(n3465), .SN(n3464), 
        .Q(iaddr[0]) );
  DFFRS_X2 ifBoi_pcOut_reg_1_ ( .D(n4708), .CK(clk), .RN(n3463), .SN(n3462), 
        .Q(iaddr[1]) );
  DFFRS_X2 ifBoi_pcOut_reg_2_ ( .D(n4703), .CK(clk), .RN(n3461), .SN(n3460), 
        .Q(iaddr[2]), .QN(n5355) );
  DFFRS_X2 ifBoi_pcOut_reg_3_ ( .D(n4698), .CK(clk), .RN(n3459), .SN(n3458), 
        .Q(iaddr[3]), .QN(n5477) );
  DFFRS_X2 ifBoi_pcOut_reg_4_ ( .D(n4693), .CK(clk), .RN(n3457), .SN(n3456), 
        .Q(iaddr[4]) );
  DFFRS_X2 ifBoi_pcOut_reg_5_ ( .D(n4688), .CK(clk), .RN(n3455), .SN(n3454), 
        .Q(iaddr[5]), .QN(n5509) );
  DFFRS_X2 ifBoi_pcOut_reg_6_ ( .D(n4683), .CK(clk), .RN(n3453), .SN(n3452), 
        .Q(iaddr[6]) );
  DFFRS_X2 ifBoi_pcOut_reg_7_ ( .D(n4678), .CK(clk), .RN(n3451), .SN(n3450), 
        .Q(iaddr[7]) );
  DFFRS_X2 ifBoi_pcOut_reg_8_ ( .D(n4673), .CK(clk), .RN(n3449), .SN(n3448), 
        .Q(iaddr[8]) );
  DFFRS_X2 ifBoi_pcOut_reg_9_ ( .D(n4668), .CK(clk), .RN(n3447), .SN(n3446), 
        .Q(iaddr[9]), .QN(n5647) );
  DFFRS_X2 ifBoi_pcOut_reg_10_ ( .D(n4663), .CK(clk), .RN(n3445), .SN(n3444), 
        .Q(iaddr[10]), .QN(n5478) );
  DFFRS_X2 ifBoi_pcOut_reg_11_ ( .D(n4658), .CK(clk), .RN(n3443), .SN(n3442), 
        .Q(iaddr[11]) );
  DFFRS_X2 ifBoi_pcOut_reg_12_ ( .D(n4653), .CK(clk), .RN(n3441), .SN(n3440), 
        .Q(iaddr[12]) );
  DFFRS_X2 ifBoi_pcOut_reg_13_ ( .D(n4648), .CK(clk), .RN(n3439), .SN(n3438), 
        .Q(iaddr[13]), .QN(n5564) );
  DFFRS_X2 ifBoi_pcOut_reg_14_ ( .D(n4643), .CK(clk), .RN(n3437), .SN(n3436), 
        .Q(iaddr[14]) );
  DFFRS_X2 ifBoi_pcOut_reg_15_ ( .D(n4638), .CK(clk), .RN(n3435), .SN(n3434), 
        .Q(iaddr[15]), .QN(n5574) );
  DFFRS_X2 ifBoi_pcOut_reg_16_ ( .D(n4633), .CK(clk), .RN(n3433), .SN(n3432), 
        .Q(iaddr[16]) );
  DFFRS_X2 ifBoi_pcOut_reg_17_ ( .D(n4628), .CK(clk), .RN(n3431), .SN(n3430), 
        .Q(iaddr[17]), .QN(n5581) );
  DFFRS_X2 ifBoi_pcOut_reg_18_ ( .D(n4623), .CK(clk), .RN(n3429), .SN(n3428), 
        .Q(iaddr[18]) );
  DFFRS_X2 ifBoi_pcOut_reg_19_ ( .D(n4618), .CK(clk), .RN(n3427), .SN(n3426), 
        .Q(iaddr[19]), .QN(n5563) );
  DFFRS_X2 ifBoi_pcOut_reg_20_ ( .D(n4613), .CK(clk), .RN(n3425), .SN(n3424), 
        .Q(iaddr[20]) );
  DFFRS_X2 ifBoi_pcOut_reg_22_ ( .D(n4603), .CK(clk), .RN(n3421), .SN(n3420), 
        .Q(iaddr[22]) );
  DFFRS_X2 ifBoi_pcOut_reg_23_ ( .D(n4598), .CK(clk), .RN(n3419), .SN(n3418), 
        .Q(iaddr[23]) );
  DFFRS_X2 ifBoi_pcOut_reg_25_ ( .D(n4588), .CK(clk), .RN(n3415), .SN(n3414), 
        .Q(iaddr[25]) );
  DFFRS_X2 ifBoi_pcOut_reg_30_ ( .D(n4563), .CK(clk), .RN(n3405), .SN(n3404), 
        .Q(iaddr[30]) );
  DFFRS_X2 ifBoi_pcOut_reg_31_ ( .D(n4558), .CK(clk), .RN(n3403), .SN(n3402), 
        .Q(iaddr[31]) );
  NAND2_X2 U2 ( .A1(regBoiz_regfile_9__9_), .A2(n6781), .ZN(n36) );
  NAND2_X2 U4 ( .A1(regBoiz_regfile_9__8_), .A2(n6780), .ZN(n38) );
  NAND2_X2 U6 ( .A1(regBoiz_regfile_9__7_), .A2(n6779), .ZN(n40) );
  NAND2_X2 U8 ( .A1(regBoiz_regfile_9__6_), .A2(n6780), .ZN(n42) );
  NAND2_X2 U10 ( .A1(regBoiz_regfile_9__5_), .A2(n6779), .ZN(n44) );
  NAND2_X2 U12 ( .A1(regBoiz_regfile_9__4_), .A2(n6779), .ZN(n46) );
  NAND2_X2 U14 ( .A1(regBoiz_regfile_9__3_), .A2(n6780), .ZN(n48) );
  NAND2_X2 U16 ( .A1(regBoiz_regfile_9__31_), .A2(n6781), .ZN(n50) );
  NAND2_X2 U18 ( .A1(regBoiz_regfile_9__30_), .A2(n6781), .ZN(n52) );
  NAND2_X2 U20 ( .A1(regBoiz_regfile_9__2_), .A2(n6781), .ZN(n54) );
  NAND2_X2 U22 ( .A1(regBoiz_regfile_9__29_), .A2(n6781), .ZN(n56) );
  NAND2_X2 U24 ( .A1(regBoiz_regfile_9__28_), .A2(n6781), .ZN(n58) );
  NAND2_X2 U26 ( .A1(regBoiz_regfile_9__27_), .A2(n6781), .ZN(n60) );
  NAND2_X2 U28 ( .A1(regBoiz_regfile_9__26_), .A2(n6781), .ZN(n62) );
  NAND2_X2 U30 ( .A1(regBoiz_regfile_9__25_), .A2(n6781), .ZN(n64) );
  NAND2_X2 U32 ( .A1(regBoiz_regfile_9__24_), .A2(n6781), .ZN(n66) );
  NAND2_X2 U34 ( .A1(regBoiz_regfile_9__23_), .A2(n6781), .ZN(n68) );
  NAND2_X2 U36 ( .A1(regBoiz_regfile_9__22_), .A2(n6781), .ZN(n70) );
  NAND2_X2 U38 ( .A1(regBoiz_regfile_9__21_), .A2(n6781), .ZN(n72) );
  NAND2_X2 U40 ( .A1(regBoiz_regfile_9__20_), .A2(n6781), .ZN(n74) );
  NAND2_X2 U42 ( .A1(regBoiz_regfile_9__1_), .A2(n6781), .ZN(n76) );
  NAND2_X2 U44 ( .A1(regBoiz_regfile_9__19_), .A2(n6781), .ZN(n78) );
  NAND2_X2 U46 ( .A1(regBoiz_regfile_9__18_), .A2(n6781), .ZN(n80) );
  NAND2_X2 U48 ( .A1(regBoiz_regfile_9__17_), .A2(n6781), .ZN(n82) );
  NAND2_X2 U50 ( .A1(regBoiz_regfile_9__16_), .A2(n6781), .ZN(n84) );
  NAND2_X2 U52 ( .A1(regBoiz_regfile_9__15_), .A2(n6780), .ZN(n86) );
  NAND2_X2 U54 ( .A1(regBoiz_regfile_9__14_), .A2(n6781), .ZN(n88) );
  NAND2_X2 U56 ( .A1(regBoiz_regfile_9__13_), .A2(n6781), .ZN(n90) );
  NAND2_X2 U58 ( .A1(regBoiz_regfile_9__12_), .A2(n6781), .ZN(n92) );
  NAND2_X2 U60 ( .A1(regBoiz_regfile_9__11_), .A2(n6781), .ZN(n94) );
  NAND2_X2 U62 ( .A1(regBoiz_regfile_9__10_), .A2(n6781), .ZN(n96) );
  NAND2_X2 U64 ( .A1(regBoiz_regfile_9__0_), .A2(n6781), .ZN(n98) );
  NAND2_X2 U65 ( .A1(n99), .A2(n100), .ZN(n34) );
  NAND2_X2 U67 ( .A1(regBoiz_regfile_8__9_), .A2(n6777), .ZN(n102) );
  NAND2_X2 U85 ( .A1(regBoiz_regfile_8__8_), .A2(n6775), .ZN(n103) );
  NAND2_X2 U87 ( .A1(regBoiz_regfile_8__7_), .A2(n6776), .ZN(n104) );
  NAND2_X2 U89 ( .A1(regBoiz_regfile_8__6_), .A2(n6775), .ZN(n105) );
  NAND2_X2 U91 ( .A1(regBoiz_regfile_8__5_), .A2(n6776), .ZN(n106) );
  NAND2_X2 U93 ( .A1(regBoiz_regfile_8__4_), .A2(n6775), .ZN(n107) );
  NAND2_X2 U95 ( .A1(regBoiz_regfile_8__3_), .A2(n6776), .ZN(n108) );
  NAND2_X2 U97 ( .A1(regBoiz_regfile_8__31_), .A2(n6775), .ZN(n109) );
  NAND2_X2 U99 ( .A1(regBoiz_regfile_8__30_), .A2(n6777), .ZN(n110) );
  NAND2_X2 U101 ( .A1(regBoiz_regfile_8__2_), .A2(n6777), .ZN(n111) );
  NAND2_X2 U103 ( .A1(regBoiz_regfile_8__29_), .A2(n6777), .ZN(n112) );
  NAND2_X2 U105 ( .A1(regBoiz_regfile_8__28_), .A2(n6777), .ZN(n113) );
  NAND2_X2 U107 ( .A1(regBoiz_regfile_8__27_), .A2(n6777), .ZN(n114) );
  NAND2_X2 U109 ( .A1(regBoiz_regfile_8__26_), .A2(n6777), .ZN(n115) );
  NAND2_X2 U111 ( .A1(regBoiz_regfile_8__25_), .A2(n6777), .ZN(n116) );
  NAND2_X2 U113 ( .A1(regBoiz_regfile_8__24_), .A2(n6777), .ZN(n117) );
  NAND2_X2 U115 ( .A1(regBoiz_regfile_8__23_), .A2(n6777), .ZN(n118) );
  NAND2_X2 U117 ( .A1(regBoiz_regfile_8__22_), .A2(n6777), .ZN(n119) );
  NAND2_X2 U119 ( .A1(regBoiz_regfile_8__21_), .A2(n6777), .ZN(n120) );
  NAND2_X2 U121 ( .A1(regBoiz_regfile_8__20_), .A2(n6777), .ZN(n121) );
  NAND2_X2 U123 ( .A1(regBoiz_regfile_8__1_), .A2(n6777), .ZN(n122) );
  NAND2_X2 U125 ( .A1(regBoiz_regfile_8__19_), .A2(n6777), .ZN(n123) );
  NAND2_X2 U127 ( .A1(regBoiz_regfile_8__18_), .A2(n6777), .ZN(n124) );
  NAND2_X2 U129 ( .A1(regBoiz_regfile_8__17_), .A2(n6777), .ZN(n125) );
  NAND2_X2 U131 ( .A1(regBoiz_regfile_8__16_), .A2(n6777), .ZN(n126) );
  NAND2_X2 U133 ( .A1(regBoiz_regfile_8__15_), .A2(n6777), .ZN(n127) );
  NAND2_X2 U135 ( .A1(regBoiz_regfile_8__14_), .A2(n6777), .ZN(n128) );
  NAND2_X2 U137 ( .A1(regBoiz_regfile_8__13_), .A2(n6777), .ZN(n129) );
  NAND2_X2 U139 ( .A1(regBoiz_regfile_8__12_), .A2(n6777), .ZN(n130) );
  NAND2_X2 U141 ( .A1(regBoiz_regfile_8__11_), .A2(n6777), .ZN(n131) );
  NAND2_X2 U143 ( .A1(regBoiz_regfile_8__10_), .A2(n6777), .ZN(n132) );
  NAND2_X2 U145 ( .A1(regBoiz_regfile_8__0_), .A2(n6777), .ZN(n133) );
  NAND2_X2 U148 ( .A1(regBoiz_regfile_7__9_), .A2(n6774), .ZN(n136) );
  NAND2_X2 U150 ( .A1(regBoiz_regfile_7__8_), .A2(n6773), .ZN(n137) );
  NAND2_X2 U156 ( .A1(regBoiz_regfile_7__5_), .A2(n6773), .ZN(n140) );
  NAND2_X2 U158 ( .A1(regBoiz_regfile_7__4_), .A2(n6772), .ZN(n141) );
  NAND2_X2 U160 ( .A1(regBoiz_regfile_7__3_), .A2(n6772), .ZN(n142) );
  NAND2_X2 U162 ( .A1(regBoiz_regfile_7__31_), .A2(n6773), .ZN(n143) );
  NAND2_X2 U164 ( .A1(regBoiz_regfile_7__30_), .A2(n6773), .ZN(n144) );
  NAND2_X2 U166 ( .A1(regBoiz_regfile_7__2_), .A2(n135), .ZN(n145) );
  NAND2_X2 U168 ( .A1(regBoiz_regfile_7__29_), .A2(n6772), .ZN(n146) );
  NAND2_X2 U170 ( .A1(regBoiz_regfile_7__28_), .A2(n135), .ZN(n147) );
  NAND2_X2 U172 ( .A1(regBoiz_regfile_7__27_), .A2(n135), .ZN(n148) );
  NAND2_X2 U174 ( .A1(regBoiz_regfile_7__26_), .A2(n135), .ZN(n149) );
  NAND2_X2 U176 ( .A1(regBoiz_regfile_7__25_), .A2(n135), .ZN(n150) );
  NAND2_X2 U178 ( .A1(regBoiz_regfile_7__24_), .A2(n135), .ZN(n151) );
  NAND2_X2 U180 ( .A1(regBoiz_regfile_7__23_), .A2(n135), .ZN(n152) );
  NAND2_X2 U182 ( .A1(regBoiz_regfile_7__22_), .A2(n135), .ZN(n153) );
  NAND2_X2 U184 ( .A1(regBoiz_regfile_7__21_), .A2(n135), .ZN(n154) );
  NAND2_X2 U186 ( .A1(regBoiz_regfile_7__20_), .A2(n135), .ZN(n155) );
  NAND2_X2 U190 ( .A1(regBoiz_regfile_7__19_), .A2(n135), .ZN(n157) );
  NAND2_X2 U192 ( .A1(regBoiz_regfile_7__18_), .A2(n6774), .ZN(n158) );
  NAND2_X2 U194 ( .A1(regBoiz_regfile_7__17_), .A2(n135), .ZN(n159) );
  NAND2_X2 U196 ( .A1(regBoiz_regfile_7__16_), .A2(n6774), .ZN(n160) );
  NAND2_X2 U198 ( .A1(regBoiz_regfile_7__15_), .A2(n6774), .ZN(n161) );
  NAND2_X2 U200 ( .A1(regBoiz_regfile_7__14_), .A2(n135), .ZN(n162) );
  NAND2_X2 U202 ( .A1(regBoiz_regfile_7__13_), .A2(n6774), .ZN(n163) );
  NAND2_X2 U204 ( .A1(regBoiz_regfile_7__12_), .A2(n6774), .ZN(n164) );
  NAND2_X2 U206 ( .A1(regBoiz_regfile_7__11_), .A2(n135), .ZN(n165) );
  NAND2_X2 U208 ( .A1(regBoiz_regfile_7__10_), .A2(n6774), .ZN(n166) );
  NAND2_X2 U210 ( .A1(regBoiz_regfile_7__0_), .A2(n135), .ZN(n167) );
  NAND2_X2 U211 ( .A1(n168), .A2(n169), .ZN(n135) );
  NAND2_X2 U213 ( .A1(regBoiz_regfile_6__9_), .A2(n6770), .ZN(n171) );
  NAND2_X2 U215 ( .A1(regBoiz_regfile_6__8_), .A2(n6769), .ZN(n172) );
  NAND2_X2 U217 ( .A1(regBoiz_regfile_6__7_), .A2(n6768), .ZN(n173) );
  NAND2_X2 U219 ( .A1(regBoiz_regfile_6__6_), .A2(n6769), .ZN(n174) );
  NAND2_X2 U221 ( .A1(regBoiz_regfile_6__5_), .A2(n6768), .ZN(n175) );
  NAND2_X2 U225 ( .A1(regBoiz_regfile_6__3_), .A2(n6769), .ZN(n177) );
  NAND2_X2 U227 ( .A1(regBoiz_regfile_6__31_), .A2(n6768), .ZN(n178) );
  NAND2_X2 U229 ( .A1(regBoiz_regfile_6__30_), .A2(n6770), .ZN(n179) );
  NAND2_X2 U231 ( .A1(regBoiz_regfile_6__2_), .A2(n6770), .ZN(n180) );
  NAND2_X2 U235 ( .A1(regBoiz_regfile_6__28_), .A2(n6770), .ZN(n182) );
  NAND2_X2 U237 ( .A1(regBoiz_regfile_6__27_), .A2(n6770), .ZN(n183) );
  NAND2_X2 U239 ( .A1(regBoiz_regfile_6__26_), .A2(n6770), .ZN(n184) );
  NAND2_X2 U241 ( .A1(regBoiz_regfile_6__25_), .A2(n6770), .ZN(n185) );
  NAND2_X2 U243 ( .A1(regBoiz_regfile_6__24_), .A2(n6770), .ZN(n186) );
  NAND2_X2 U245 ( .A1(regBoiz_regfile_6__23_), .A2(n6770), .ZN(n187) );
  NAND2_X2 U247 ( .A1(regBoiz_regfile_6__22_), .A2(n6770), .ZN(n188) );
  NAND2_X2 U249 ( .A1(regBoiz_regfile_6__21_), .A2(n6770), .ZN(n189) );
  NAND2_X2 U251 ( .A1(regBoiz_regfile_6__20_), .A2(n6770), .ZN(n190) );
  NAND2_X2 U253 ( .A1(regBoiz_regfile_6__1_), .A2(n6770), .ZN(n191) );
  NAND2_X2 U255 ( .A1(regBoiz_regfile_6__19_), .A2(n6770), .ZN(n192) );
  NAND2_X2 U257 ( .A1(regBoiz_regfile_6__18_), .A2(n6770), .ZN(n193) );
  NAND2_X2 U259 ( .A1(regBoiz_regfile_6__17_), .A2(n6770), .ZN(n194) );
  NAND2_X2 U261 ( .A1(regBoiz_regfile_6__16_), .A2(n6770), .ZN(n195) );
  NAND2_X2 U263 ( .A1(regBoiz_regfile_6__15_), .A2(n6770), .ZN(n196) );
  NAND2_X2 U265 ( .A1(regBoiz_regfile_6__14_), .A2(n6770), .ZN(n197) );
  NAND2_X2 U267 ( .A1(regBoiz_regfile_6__13_), .A2(n6770), .ZN(n198) );
  NAND2_X2 U269 ( .A1(regBoiz_regfile_6__12_), .A2(n6770), .ZN(n199) );
  NAND2_X2 U271 ( .A1(regBoiz_regfile_6__11_), .A2(n6770), .ZN(n200) );
  NAND2_X2 U273 ( .A1(regBoiz_regfile_6__10_), .A2(n6770), .ZN(n201) );
  NAND2_X2 U275 ( .A1(regBoiz_regfile_6__0_), .A2(n6770), .ZN(n202) );
  NAND2_X2 U278 ( .A1(regBoiz_regfile_5__9_), .A2(n6767), .ZN(n205) );
  NAND2_X2 U280 ( .A1(regBoiz_regfile_5__8_), .A2(n6765), .ZN(n206) );
  NAND2_X2 U282 ( .A1(regBoiz_regfile_5__7_), .A2(n6766), .ZN(n207) );
  NAND2_X2 U284 ( .A1(regBoiz_regfile_5__6_), .A2(n6765), .ZN(n208) );
  NAND2_X2 U286 ( .A1(regBoiz_regfile_5__5_), .A2(n6766), .ZN(n209) );
  NAND2_X2 U288 ( .A1(regBoiz_regfile_5__4_), .A2(n6766), .ZN(n210) );
  NAND2_X2 U290 ( .A1(regBoiz_regfile_5__3_), .A2(n6765), .ZN(n211) );
  NAND2_X2 U292 ( .A1(regBoiz_regfile_5__31_), .A2(n6765), .ZN(n212) );
  NAND2_X2 U294 ( .A1(regBoiz_regfile_5__30_), .A2(n6767), .ZN(n213) );
  NAND2_X2 U296 ( .A1(regBoiz_regfile_5__2_), .A2(n6767), .ZN(n214) );
  NAND2_X2 U298 ( .A1(regBoiz_regfile_5__29_), .A2(n6767), .ZN(n215) );
  NAND2_X2 U300 ( .A1(regBoiz_regfile_5__28_), .A2(n6767), .ZN(n216) );
  NAND2_X2 U302 ( .A1(regBoiz_regfile_5__27_), .A2(n6767), .ZN(n217) );
  NAND2_X2 U304 ( .A1(regBoiz_regfile_5__26_), .A2(n6767), .ZN(n218) );
  NAND2_X2 U306 ( .A1(regBoiz_regfile_5__25_), .A2(n6767), .ZN(n219) );
  NAND2_X2 U308 ( .A1(regBoiz_regfile_5__24_), .A2(n6767), .ZN(n220) );
  NAND2_X2 U310 ( .A1(regBoiz_regfile_5__23_), .A2(n6767), .ZN(n221) );
  NAND2_X2 U312 ( .A1(regBoiz_regfile_5__22_), .A2(n6767), .ZN(n222) );
  NAND2_X2 U314 ( .A1(regBoiz_regfile_5__21_), .A2(n6767), .ZN(n223) );
  NAND2_X2 U316 ( .A1(regBoiz_regfile_5__20_), .A2(n6767), .ZN(n224) );
  NAND2_X2 U318 ( .A1(regBoiz_regfile_5__1_), .A2(n6767), .ZN(n225) );
  NAND2_X2 U320 ( .A1(regBoiz_regfile_5__19_), .A2(n6767), .ZN(n226) );
  NAND2_X2 U322 ( .A1(regBoiz_regfile_5__18_), .A2(n6767), .ZN(n227) );
  NAND2_X2 U324 ( .A1(regBoiz_regfile_5__17_), .A2(n6767), .ZN(n228) );
  NAND2_X2 U326 ( .A1(regBoiz_regfile_5__16_), .A2(n6767), .ZN(n229) );
  NAND2_X2 U328 ( .A1(regBoiz_regfile_5__15_), .A2(n6767), .ZN(n230) );
  NAND2_X2 U330 ( .A1(regBoiz_regfile_5__14_), .A2(n6767), .ZN(n231) );
  NAND2_X2 U332 ( .A1(regBoiz_regfile_5__13_), .A2(n6767), .ZN(n232) );
  NAND2_X2 U334 ( .A1(regBoiz_regfile_5__12_), .A2(n6767), .ZN(n233) );
  NAND2_X2 U336 ( .A1(regBoiz_regfile_5__11_), .A2(n6767), .ZN(n234) );
  NAND2_X2 U338 ( .A1(regBoiz_regfile_5__10_), .A2(n6767), .ZN(n235) );
  NAND2_X2 U340 ( .A1(regBoiz_regfile_5__0_), .A2(n6767), .ZN(n236) );
  NAND2_X2 U343 ( .A1(regBoiz_regfile_4__9_), .A2(n6762), .ZN(n238) );
  NAND2_X2 U345 ( .A1(regBoiz_regfile_4__8_), .A2(n6761), .ZN(n239) );
  NAND2_X2 U347 ( .A1(regBoiz_regfile_4__7_), .A2(n6762), .ZN(n240) );
  NAND2_X2 U349 ( .A1(regBoiz_regfile_4__6_), .A2(n6761), .ZN(n241) );
  NAND2_X2 U351 ( .A1(regBoiz_regfile_4__5_), .A2(n6762), .ZN(n242) );
  NAND2_X2 U353 ( .A1(regBoiz_regfile_4__4_), .A2(n6761), .ZN(n243) );
  NAND2_X2 U355 ( .A1(regBoiz_regfile_4__3_), .A2(n6762), .ZN(n244) );
  NAND2_X2 U357 ( .A1(regBoiz_regfile_4__31_), .A2(n6763), .ZN(n245) );
  NAND2_X2 U359 ( .A1(regBoiz_regfile_4__30_), .A2(n6763), .ZN(n246) );
  NAND2_X2 U361 ( .A1(regBoiz_regfile_4__2_), .A2(n6763), .ZN(n247) );
  NAND2_X2 U363 ( .A1(regBoiz_regfile_4__29_), .A2(n6763), .ZN(n248) );
  NAND2_X2 U365 ( .A1(regBoiz_regfile_4__28_), .A2(n6763), .ZN(n249) );
  NAND2_X2 U367 ( .A1(regBoiz_regfile_4__27_), .A2(n6763), .ZN(n250) );
  NAND2_X2 U369 ( .A1(regBoiz_regfile_4__26_), .A2(n6763), .ZN(n251) );
  NAND2_X2 U371 ( .A1(regBoiz_regfile_4__25_), .A2(n6763), .ZN(n252) );
  NAND2_X2 U373 ( .A1(regBoiz_regfile_4__24_), .A2(n6763), .ZN(n253) );
  NAND2_X2 U375 ( .A1(regBoiz_regfile_4__23_), .A2(n6763), .ZN(n254) );
  NAND2_X2 U377 ( .A1(regBoiz_regfile_4__22_), .A2(n6763), .ZN(n255) );
  NAND2_X2 U379 ( .A1(regBoiz_regfile_4__21_), .A2(n6763), .ZN(n256) );
  NAND2_X2 U381 ( .A1(regBoiz_regfile_4__20_), .A2(n6763), .ZN(n257) );
  NAND2_X2 U383 ( .A1(regBoiz_regfile_4__1_), .A2(n6763), .ZN(n258) );
  NAND2_X2 U385 ( .A1(regBoiz_regfile_4__19_), .A2(n6763), .ZN(n259) );
  NAND2_X2 U387 ( .A1(regBoiz_regfile_4__18_), .A2(n6763), .ZN(n260) );
  NAND2_X2 U389 ( .A1(regBoiz_regfile_4__17_), .A2(n6763), .ZN(n261) );
  NAND2_X2 U391 ( .A1(regBoiz_regfile_4__16_), .A2(n6761), .ZN(n262) );
  NAND2_X2 U393 ( .A1(regBoiz_regfile_4__15_), .A2(n6763), .ZN(n263) );
  NAND2_X2 U395 ( .A1(regBoiz_regfile_4__14_), .A2(n6763), .ZN(n264) );
  NAND2_X2 U397 ( .A1(regBoiz_regfile_4__13_), .A2(n6762), .ZN(n265) );
  NAND2_X2 U399 ( .A1(regBoiz_regfile_4__12_), .A2(n6763), .ZN(n266) );
  NAND2_X2 U401 ( .A1(regBoiz_regfile_4__11_), .A2(n6763), .ZN(n267) );
  NAND2_X2 U403 ( .A1(regBoiz_regfile_4__10_), .A2(n6763), .ZN(n268) );
  NAND2_X2 U405 ( .A1(regBoiz_regfile_4__0_), .A2(n6763), .ZN(n269) );
  NAND2_X2 U406 ( .A1(n169), .A2(n134), .ZN(n237) );
  AND2_X2 U407 ( .A1(n270), .A2(n271), .ZN(n169) );
  NAND2_X2 U409 ( .A1(regBoiz_regfile_3__9_), .A2(n6760), .ZN(n273) );
  NAND2_X2 U411 ( .A1(regBoiz_regfile_3__8_), .A2(n6758), .ZN(n274) );
  NAND2_X2 U413 ( .A1(regBoiz_regfile_3__7_), .A2(n6759), .ZN(n275) );
  NAND2_X2 U415 ( .A1(regBoiz_regfile_3__6_), .A2(n6758), .ZN(n276) );
  NAND2_X2 U417 ( .A1(regBoiz_regfile_3__5_), .A2(n6759), .ZN(n277) );
  NAND2_X2 U421 ( .A1(regBoiz_regfile_3__3_), .A2(n6758), .ZN(n279) );
  NAND2_X2 U423 ( .A1(regBoiz_regfile_3__31_), .A2(n6759), .ZN(n280) );
  NAND2_X2 U425 ( .A1(regBoiz_regfile_3__30_), .A2(n6760), .ZN(n281) );
  NAND2_X2 U427 ( .A1(regBoiz_regfile_3__2_), .A2(n6760), .ZN(n282) );
  NAND2_X2 U429 ( .A1(regBoiz_regfile_3__29_), .A2(n6760), .ZN(n283) );
  NAND2_X2 U431 ( .A1(regBoiz_regfile_3__28_), .A2(n6760), .ZN(n284) );
  NAND2_X2 U433 ( .A1(regBoiz_regfile_3__27_), .A2(n6760), .ZN(n285) );
  NAND2_X2 U435 ( .A1(regBoiz_regfile_3__26_), .A2(n6760), .ZN(n286) );
  NAND2_X2 U437 ( .A1(regBoiz_regfile_3__25_), .A2(n6760), .ZN(n287) );
  NAND2_X2 U439 ( .A1(regBoiz_regfile_3__24_), .A2(n6760), .ZN(n288) );
  NAND2_X2 U441 ( .A1(regBoiz_regfile_3__23_), .A2(n6760), .ZN(n289) );
  NAND2_X2 U443 ( .A1(regBoiz_regfile_3__22_), .A2(n6760), .ZN(n290) );
  NAND2_X2 U445 ( .A1(regBoiz_regfile_3__21_), .A2(n6760), .ZN(n291) );
  NAND2_X2 U447 ( .A1(regBoiz_regfile_3__20_), .A2(n6760), .ZN(n292) );
  NAND2_X2 U449 ( .A1(regBoiz_regfile_3__1_), .A2(n6760), .ZN(n293) );
  NAND2_X2 U451 ( .A1(regBoiz_regfile_3__19_), .A2(n6760), .ZN(n294) );
  NAND2_X2 U453 ( .A1(regBoiz_regfile_3__18_), .A2(n6760), .ZN(n295) );
  NAND2_X2 U455 ( .A1(regBoiz_regfile_3__17_), .A2(n6760), .ZN(n296) );
  NAND2_X2 U457 ( .A1(regBoiz_regfile_3__16_), .A2(n6760), .ZN(n297) );
  NAND2_X2 U459 ( .A1(regBoiz_regfile_3__15_), .A2(n6760), .ZN(n298) );
  NAND2_X2 U461 ( .A1(regBoiz_regfile_3__14_), .A2(n6760), .ZN(n299) );
  NAND2_X2 U463 ( .A1(regBoiz_regfile_3__13_), .A2(n6760), .ZN(n300) );
  NAND2_X2 U465 ( .A1(regBoiz_regfile_3__12_), .A2(n6760), .ZN(n301) );
  NAND2_X2 U467 ( .A1(regBoiz_regfile_3__11_), .A2(n6760), .ZN(n302) );
  NAND2_X2 U469 ( .A1(regBoiz_regfile_3__10_), .A2(n6760), .ZN(n303) );
  NAND2_X2 U471 ( .A1(regBoiz_regfile_3__0_), .A2(n6760), .ZN(n304) );
  NAND2_X2 U474 ( .A1(regBoiz_regfile_31__9_), .A2(n6757), .ZN(n307) );
  NAND2_X2 U476 ( .A1(regBoiz_regfile_31__8_), .A2(n6756), .ZN(n308) );
  NAND2_X2 U478 ( .A1(regBoiz_regfile_31__7_), .A2(n6756), .ZN(n309) );
  NAND2_X2 U482 ( .A1(regBoiz_regfile_31__5_), .A2(n6756), .ZN(n311) );
  NAND2_X2 U484 ( .A1(regBoiz_regfile_31__4_), .A2(n6756), .ZN(n312) );
  NAND2_X2 U486 ( .A1(regBoiz_regfile_31__3_), .A2(n6756), .ZN(n313) );
  NAND2_X2 U488 ( .A1(regBoiz_regfile_31__31_), .A2(n6756), .ZN(n314) );
  NAND2_X2 U490 ( .A1(regBoiz_regfile_31__30_), .A2(n6757), .ZN(n315) );
  NAND2_X2 U496 ( .A1(regBoiz_regfile_31__28_), .A2(n6757), .ZN(n318) );
  NAND2_X2 U498 ( .A1(regBoiz_regfile_31__27_), .A2(n6757), .ZN(n319) );
  NAND2_X2 U500 ( .A1(regBoiz_regfile_31__26_), .A2(n6757), .ZN(n320) );
  NAND2_X2 U502 ( .A1(regBoiz_regfile_31__25_), .A2(n6757), .ZN(n321) );
  NAND2_X2 U504 ( .A1(regBoiz_regfile_31__24_), .A2(n6757), .ZN(n322) );
  NAND2_X2 U506 ( .A1(regBoiz_regfile_31__23_), .A2(n6757), .ZN(n323) );
  NAND2_X2 U508 ( .A1(regBoiz_regfile_31__22_), .A2(n6757), .ZN(n324) );
  NAND2_X2 U510 ( .A1(regBoiz_regfile_31__21_), .A2(n6757), .ZN(n325) );
  NAND2_X2 U512 ( .A1(regBoiz_regfile_31__20_), .A2(n6757), .ZN(n326) );
  NAND2_X2 U516 ( .A1(regBoiz_regfile_31__19_), .A2(n6757), .ZN(n328) );
  NAND2_X2 U518 ( .A1(regBoiz_regfile_31__18_), .A2(n6757), .ZN(n329) );
  NAND2_X2 U520 ( .A1(regBoiz_regfile_31__17_), .A2(n6757), .ZN(n330) );
  NAND2_X2 U522 ( .A1(regBoiz_regfile_31__16_), .A2(n6757), .ZN(n331) );
  NAND2_X2 U524 ( .A1(regBoiz_regfile_31__15_), .A2(n6757), .ZN(n332) );
  NAND2_X2 U526 ( .A1(regBoiz_regfile_31__14_), .A2(n6757), .ZN(n333) );
  NAND2_X2 U532 ( .A1(regBoiz_regfile_31__11_), .A2(n6757), .ZN(n336) );
  NAND2_X2 U536 ( .A1(regBoiz_regfile_31__0_), .A2(n6757), .ZN(n338) );
  NAND2_X2 U539 ( .A1(regBoiz_regfile_30__9_), .A2(n340), .ZN(n341) );
  NAND2_X2 U541 ( .A1(regBoiz_regfile_30__8_), .A2(n6753), .ZN(n342) );
  NAND2_X2 U543 ( .A1(regBoiz_regfile_30__7_), .A2(n6752), .ZN(n343) );
  NAND2_X2 U545 ( .A1(regBoiz_regfile_30__6_), .A2(n6753), .ZN(n344) );
  NAND2_X2 U549 ( .A1(regBoiz_regfile_30__4_), .A2(n6753), .ZN(n346) );
  NAND2_X2 U551 ( .A1(regBoiz_regfile_30__3_), .A2(n6752), .ZN(n347) );
  NAND2_X2 U553 ( .A1(regBoiz_regfile_30__31_), .A2(n6752), .ZN(n348) );
  NAND2_X2 U555 ( .A1(regBoiz_regfile_30__30_), .A2(n340), .ZN(n349) );
  NAND2_X2 U557 ( .A1(regBoiz_regfile_30__2_), .A2(n340), .ZN(n350) );
  NAND2_X2 U561 ( .A1(regBoiz_regfile_30__28_), .A2(n340), .ZN(n352) );
  NAND2_X2 U563 ( .A1(regBoiz_regfile_30__27_), .A2(n340), .ZN(n353) );
  NAND2_X2 U565 ( .A1(regBoiz_regfile_30__26_), .A2(n340), .ZN(n354) );
  NAND2_X2 U567 ( .A1(regBoiz_regfile_30__25_), .A2(n340), .ZN(n355) );
  NAND2_X2 U569 ( .A1(regBoiz_regfile_30__24_), .A2(n340), .ZN(n356) );
  NAND2_X2 U571 ( .A1(regBoiz_regfile_30__23_), .A2(n340), .ZN(n357) );
  NAND2_X2 U573 ( .A1(regBoiz_regfile_30__22_), .A2(n340), .ZN(n358) );
  NAND2_X2 U575 ( .A1(regBoiz_regfile_30__21_), .A2(n340), .ZN(n359) );
  NAND2_X2 U577 ( .A1(regBoiz_regfile_30__20_), .A2(n340), .ZN(n360) );
  NAND2_X2 U579 ( .A1(regBoiz_regfile_30__1_), .A2(n340), .ZN(n361) );
  NAND2_X2 U581 ( .A1(regBoiz_regfile_30__19_), .A2(n340), .ZN(n362) );
  NAND2_X2 U583 ( .A1(regBoiz_regfile_30__18_), .A2(n340), .ZN(n363) );
  NAND2_X2 U585 ( .A1(regBoiz_regfile_30__17_), .A2(n340), .ZN(n364) );
  NAND2_X2 U587 ( .A1(regBoiz_regfile_30__16_), .A2(n340), .ZN(n365) );
  NAND2_X2 U589 ( .A1(regBoiz_regfile_30__15_), .A2(n340), .ZN(n366) );
  NAND2_X2 U591 ( .A1(regBoiz_regfile_30__14_), .A2(n340), .ZN(n367) );
  NAND2_X2 U593 ( .A1(regBoiz_regfile_30__13_), .A2(n340), .ZN(n368) );
  NAND2_X2 U595 ( .A1(regBoiz_regfile_30__12_), .A2(n340), .ZN(n369) );
  NAND2_X2 U597 ( .A1(regBoiz_regfile_30__11_), .A2(n340), .ZN(n370) );
  NAND2_X2 U599 ( .A1(regBoiz_regfile_30__10_), .A2(n340), .ZN(n371) );
  NAND2_X2 U601 ( .A1(regBoiz_regfile_30__0_), .A2(n340), .ZN(n372) );
  NAND2_X2 U602 ( .A1(n339), .A2(n203), .ZN(n340) );
  NAND2_X2 U604 ( .A1(regBoiz_regfile_2__9_), .A2(net367221), .ZN(n374) );
  NAND2_X2 U606 ( .A1(regBoiz_regfile_2__8_), .A2(net367217), .ZN(n375) );
  NAND2_X2 U608 ( .A1(regBoiz_regfile_2__7_), .A2(net367217), .ZN(n376) );
  NAND2_X2 U610 ( .A1(regBoiz_regfile_2__6_), .A2(net367215), .ZN(n377) );
  NAND2_X2 U612 ( .A1(regBoiz_regfile_2__5_), .A2(net367217), .ZN(n378) );
  NAND2_X2 U614 ( .A1(regBoiz_regfile_2__4_), .A2(net367215), .ZN(n379) );
  NAND2_X2 U616 ( .A1(regBoiz_regfile_2__3_), .A2(net367221), .ZN(n380) );
  NAND2_X2 U618 ( .A1(regBoiz_regfile_2__31_), .A2(net367215), .ZN(n381) );
  NAND2_X2 U620 ( .A1(regBoiz_regfile_2__30_), .A2(net367221), .ZN(n382) );
  NAND2_X2 U622 ( .A1(regBoiz_regfile_2__2_), .A2(net367221), .ZN(n383) );
  NAND2_X2 U624 ( .A1(regBoiz_regfile_2__29_), .A2(net367221), .ZN(n384) );
  NAND2_X2 U626 ( .A1(regBoiz_regfile_2__28_), .A2(net367221), .ZN(n385) );
  NAND2_X2 U630 ( .A1(regBoiz_regfile_2__26_), .A2(net367221), .ZN(n387) );
  NAND2_X2 U632 ( .A1(regBoiz_regfile_2__25_), .A2(net367221), .ZN(n388) );
  NAND2_X2 U634 ( .A1(regBoiz_regfile_2__24_), .A2(net367221), .ZN(n389) );
  NAND2_X2 U636 ( .A1(regBoiz_regfile_2__23_), .A2(net367221), .ZN(n390) );
  NAND2_X2 U638 ( .A1(regBoiz_regfile_2__22_), .A2(net367221), .ZN(n391) );
  NAND2_X2 U640 ( .A1(regBoiz_regfile_2__21_), .A2(net367221), .ZN(n392) );
  NAND2_X2 U642 ( .A1(regBoiz_regfile_2__20_), .A2(net367221), .ZN(n393) );
  NAND2_X2 U644 ( .A1(regBoiz_regfile_2__1_), .A2(net367221), .ZN(n394) );
  NAND2_X2 U646 ( .A1(regBoiz_regfile_2__19_), .A2(net367221), .ZN(n395) );
  NAND2_X2 U648 ( .A1(regBoiz_regfile_2__18_), .A2(net367221), .ZN(n396) );
  NAND2_X2 U650 ( .A1(regBoiz_regfile_2__17_), .A2(net367221), .ZN(n397) );
  NAND2_X2 U652 ( .A1(regBoiz_regfile_2__16_), .A2(net367215), .ZN(n398) );
  NAND2_X2 U654 ( .A1(regBoiz_regfile_2__15_), .A2(net367221), .ZN(n399) );
  NAND2_X2 U656 ( .A1(regBoiz_regfile_2__14_), .A2(net367221), .ZN(n400) );
  NAND2_X2 U658 ( .A1(regBoiz_regfile_2__13_), .A2(net367217), .ZN(n401) );
  NAND2_X2 U660 ( .A1(regBoiz_regfile_2__12_), .A2(net367221), .ZN(n402) );
  NAND2_X2 U662 ( .A1(regBoiz_regfile_2__11_), .A2(net367221), .ZN(n403) );
  NAND2_X2 U664 ( .A1(regBoiz_regfile_2__10_), .A2(net367221), .ZN(n404) );
  NAND2_X2 U666 ( .A1(regBoiz_regfile_2__0_), .A2(net367221), .ZN(n405) );
  NAND2_X2 U667 ( .A1(n305), .A2(n203), .ZN(n373) );
  NAND2_X2 U669 ( .A1(regBoiz_regfile_29__9_), .A2(n6751), .ZN(n407) );
  NAND2_X2 U671 ( .A1(regBoiz_regfile_29__8_), .A2(n6750), .ZN(n408) );
  NAND2_X2 U673 ( .A1(regBoiz_regfile_29__7_), .A2(n6749), .ZN(n409) );
  NAND2_X2 U675 ( .A1(regBoiz_regfile_29__6_), .A2(n6750), .ZN(n410) );
  NAND2_X2 U677 ( .A1(regBoiz_regfile_29__5_), .A2(n6749), .ZN(n411) );
  NAND2_X2 U679 ( .A1(regBoiz_regfile_29__4_), .A2(n6750), .ZN(n412) );
  NAND2_X2 U681 ( .A1(regBoiz_regfile_29__3_), .A2(n6749), .ZN(n413) );
  NAND2_X2 U683 ( .A1(regBoiz_regfile_29__31_), .A2(n6749), .ZN(n414) );
  NAND2_X2 U685 ( .A1(regBoiz_regfile_29__30_), .A2(n6751), .ZN(n415) );
  NAND2_X2 U687 ( .A1(regBoiz_regfile_29__2_), .A2(n6751), .ZN(n416) );
  NAND2_X2 U689 ( .A1(regBoiz_regfile_29__29_), .A2(n6751), .ZN(n417) );
  NAND2_X2 U691 ( .A1(regBoiz_regfile_29__28_), .A2(n6751), .ZN(n418) );
  NAND2_X2 U693 ( .A1(regBoiz_regfile_29__27_), .A2(n6751), .ZN(n419) );
  NAND2_X2 U695 ( .A1(regBoiz_regfile_29__26_), .A2(n6751), .ZN(n420) );
  NAND2_X2 U697 ( .A1(regBoiz_regfile_29__25_), .A2(n6751), .ZN(n421) );
  NAND2_X2 U699 ( .A1(regBoiz_regfile_29__24_), .A2(n6751), .ZN(n422) );
  NAND2_X2 U703 ( .A1(regBoiz_regfile_29__22_), .A2(n6751), .ZN(n424) );
  NAND2_X2 U705 ( .A1(regBoiz_regfile_29__21_), .A2(n6751), .ZN(n425) );
  NAND2_X2 U707 ( .A1(regBoiz_regfile_29__20_), .A2(n6751), .ZN(n426) );
  NAND2_X2 U711 ( .A1(regBoiz_regfile_29__19_), .A2(n6751), .ZN(n428) );
  NAND2_X2 U713 ( .A1(regBoiz_regfile_29__18_), .A2(n6751), .ZN(n429) );
  NAND2_X2 U715 ( .A1(regBoiz_regfile_29__17_), .A2(n6751), .ZN(n430) );
  NAND2_X2 U717 ( .A1(regBoiz_regfile_29__16_), .A2(n6751), .ZN(n431) );
  NAND2_X2 U719 ( .A1(regBoiz_regfile_29__15_), .A2(n6751), .ZN(n432) );
  NAND2_X2 U721 ( .A1(regBoiz_regfile_29__14_), .A2(n6751), .ZN(n433) );
  NAND2_X2 U723 ( .A1(regBoiz_regfile_29__13_), .A2(n6751), .ZN(n434) );
  NAND2_X2 U725 ( .A1(regBoiz_regfile_29__12_), .A2(n6751), .ZN(n435) );
  NAND2_X2 U727 ( .A1(regBoiz_regfile_29__11_), .A2(n6751), .ZN(n436) );
  NAND2_X2 U731 ( .A1(regBoiz_regfile_29__0_), .A2(n6751), .ZN(n438) );
  NAND2_X2 U736 ( .A1(regBoiz_regfile_28__8_), .A2(n6747), .ZN(n441) );
  NAND2_X2 U738 ( .A1(regBoiz_regfile_28__7_), .A2(n6747), .ZN(n442) );
  NAND2_X2 U740 ( .A1(regBoiz_regfile_28__6_), .A2(n6747), .ZN(n443) );
  NAND2_X2 U742 ( .A1(regBoiz_regfile_28__5_), .A2(n6747), .ZN(n444) );
  NAND2_X2 U746 ( .A1(regBoiz_regfile_28__3_), .A2(n6747), .ZN(n446) );
  NAND2_X2 U748 ( .A1(regBoiz_regfile_28__31_), .A2(n6748), .ZN(n447) );
  NAND2_X2 U750 ( .A1(regBoiz_regfile_28__30_), .A2(n6748), .ZN(n448) );
  NAND2_X2 U752 ( .A1(regBoiz_regfile_28__2_), .A2(n6748), .ZN(n449) );
  NAND2_X2 U754 ( .A1(regBoiz_regfile_28__29_), .A2(n6748), .ZN(n450) );
  NAND2_X2 U756 ( .A1(regBoiz_regfile_28__28_), .A2(n6748), .ZN(n451) );
  NAND2_X2 U758 ( .A1(regBoiz_regfile_28__27_), .A2(n6748), .ZN(n452) );
  NAND2_X2 U760 ( .A1(regBoiz_regfile_28__26_), .A2(n6748), .ZN(n453) );
  NAND2_X2 U762 ( .A1(regBoiz_regfile_28__25_), .A2(n6748), .ZN(n454) );
  NAND2_X2 U764 ( .A1(regBoiz_regfile_28__24_), .A2(n6748), .ZN(n455) );
  NAND2_X2 U766 ( .A1(regBoiz_regfile_28__23_), .A2(n6748), .ZN(n456) );
  NAND2_X2 U768 ( .A1(regBoiz_regfile_28__22_), .A2(n6748), .ZN(n457) );
  NAND2_X2 U770 ( .A1(regBoiz_regfile_28__21_), .A2(n6748), .ZN(n458) );
  NAND2_X2 U772 ( .A1(regBoiz_regfile_28__20_), .A2(n6748), .ZN(n459) );
  NAND2_X2 U774 ( .A1(regBoiz_regfile_28__1_), .A2(n6748), .ZN(n460) );
  NAND2_X2 U776 ( .A1(regBoiz_regfile_28__19_), .A2(n6748), .ZN(n461) );
  NAND2_X2 U778 ( .A1(regBoiz_regfile_28__18_), .A2(n6748), .ZN(n462) );
  NAND2_X2 U780 ( .A1(regBoiz_regfile_28__17_), .A2(n6748), .ZN(n463) );
  NAND2_X2 U782 ( .A1(regBoiz_regfile_28__16_), .A2(n6747), .ZN(n464) );
  NAND2_X2 U784 ( .A1(regBoiz_regfile_28__15_), .A2(n6748), .ZN(n465) );
  NAND2_X2 U786 ( .A1(regBoiz_regfile_28__14_), .A2(n6748), .ZN(n466) );
  NAND2_X2 U788 ( .A1(regBoiz_regfile_28__13_), .A2(n6747), .ZN(n467) );
  NAND2_X2 U790 ( .A1(regBoiz_regfile_28__12_), .A2(n6748), .ZN(n468) );
  NAND2_X2 U792 ( .A1(regBoiz_regfile_28__11_), .A2(n6748), .ZN(n469) );
  NAND2_X2 U796 ( .A1(regBoiz_regfile_28__0_), .A2(n6748), .ZN(n471) );
  NAND2_X2 U797 ( .A1(n339), .A2(n134), .ZN(n439) );
  AND2_X2 U798 ( .A1(n472), .A2(wbRwh[2]), .ZN(n339) );
  NAND2_X2 U800 ( .A1(regBoiz_regfile_27__9_), .A2(n6745), .ZN(n474) );
  NAND2_X2 U802 ( .A1(regBoiz_regfile_27__8_), .A2(n6743), .ZN(n475) );
  NAND2_X2 U804 ( .A1(regBoiz_regfile_27__7_), .A2(n6744), .ZN(n476) );
  NAND2_X2 U808 ( .A1(regBoiz_regfile_27__5_), .A2(n6744), .ZN(n478) );
  NAND2_X2 U810 ( .A1(regBoiz_regfile_27__4_), .A2(n6743), .ZN(n479) );
  NAND2_X2 U812 ( .A1(regBoiz_regfile_27__3_), .A2(n6744), .ZN(n480) );
  NAND2_X2 U814 ( .A1(regBoiz_regfile_27__31_), .A2(n6743), .ZN(n481) );
  NAND2_X2 U816 ( .A1(regBoiz_regfile_27__30_), .A2(n6745), .ZN(n482) );
  NAND2_X2 U818 ( .A1(regBoiz_regfile_27__2_), .A2(n6745), .ZN(n483) );
  NAND2_X2 U820 ( .A1(regBoiz_regfile_27__29_), .A2(n6745), .ZN(n484) );
  NAND2_X2 U822 ( .A1(regBoiz_regfile_27__28_), .A2(n6745), .ZN(n485) );
  NAND2_X2 U824 ( .A1(regBoiz_regfile_27__27_), .A2(n6745), .ZN(n486) );
  NAND2_X2 U826 ( .A1(regBoiz_regfile_27__26_), .A2(n6745), .ZN(n487) );
  NAND2_X2 U828 ( .A1(regBoiz_regfile_27__25_), .A2(n6745), .ZN(n488) );
  NAND2_X2 U830 ( .A1(regBoiz_regfile_27__24_), .A2(n6745), .ZN(n489) );
  NAND2_X2 U834 ( .A1(regBoiz_regfile_27__22_), .A2(n6745), .ZN(n491) );
  NAND2_X2 U836 ( .A1(regBoiz_regfile_27__21_), .A2(n6745), .ZN(n492) );
  NAND2_X2 U838 ( .A1(regBoiz_regfile_27__20_), .A2(n6745), .ZN(n493) );
  NAND2_X2 U842 ( .A1(regBoiz_regfile_27__19_), .A2(n6745), .ZN(n495) );
  NAND2_X2 U848 ( .A1(regBoiz_regfile_27__16_), .A2(n6745), .ZN(n498) );
  NAND2_X2 U850 ( .A1(regBoiz_regfile_27__15_), .A2(n6745), .ZN(n499) );
  NAND2_X2 U852 ( .A1(regBoiz_regfile_27__14_), .A2(n6745), .ZN(n500) );
  NAND2_X2 U854 ( .A1(regBoiz_regfile_27__13_), .A2(n6745), .ZN(n501) );
  NAND2_X2 U856 ( .A1(regBoiz_regfile_27__12_), .A2(n6745), .ZN(n502) );
  NAND2_X2 U858 ( .A1(regBoiz_regfile_27__11_), .A2(n6745), .ZN(n503) );
  NAND2_X2 U862 ( .A1(regBoiz_regfile_27__0_), .A2(n6745), .ZN(n505) );
  NAND2_X2 U865 ( .A1(regBoiz_regfile_26__9_), .A2(n6740), .ZN(n508) );
  NAND2_X2 U867 ( .A1(regBoiz_regfile_26__8_), .A2(n6740), .ZN(n509) );
  NAND2_X2 U869 ( .A1(regBoiz_regfile_26__7_), .A2(n6741), .ZN(n510) );
  NAND2_X2 U871 ( .A1(regBoiz_regfile_26__6_), .A2(n6740), .ZN(n511) );
  NAND2_X2 U873 ( .A1(regBoiz_regfile_26__5_), .A2(n6741), .ZN(n512) );
  NAND2_X2 U877 ( .A1(regBoiz_regfile_26__3_), .A2(n6740), .ZN(n514) );
  NAND2_X2 U879 ( .A1(regBoiz_regfile_26__31_), .A2(n6741), .ZN(n515) );
  NAND2_X2 U881 ( .A1(regBoiz_regfile_26__30_), .A2(n6742), .ZN(n516) );
  NAND2_X2 U883 ( .A1(regBoiz_regfile_26__2_), .A2(n6742), .ZN(n517) );
  NAND2_X2 U885 ( .A1(regBoiz_regfile_26__29_), .A2(n6742), .ZN(n518) );
  NAND2_X2 U887 ( .A1(regBoiz_regfile_26__28_), .A2(n6742), .ZN(n519) );
  NAND2_X2 U889 ( .A1(regBoiz_regfile_26__27_), .A2(n6742), .ZN(n520) );
  NAND2_X2 U891 ( .A1(regBoiz_regfile_26__26_), .A2(n6742), .ZN(n521) );
  NAND2_X2 U893 ( .A1(regBoiz_regfile_26__25_), .A2(n6742), .ZN(n522) );
  NAND2_X2 U895 ( .A1(regBoiz_regfile_26__24_), .A2(n6742), .ZN(n523) );
  NAND2_X2 U897 ( .A1(regBoiz_regfile_26__23_), .A2(n6742), .ZN(n524) );
  NAND2_X2 U899 ( .A1(regBoiz_regfile_26__22_), .A2(n6742), .ZN(n525) );
  NAND2_X2 U901 ( .A1(regBoiz_regfile_26__21_), .A2(n6742), .ZN(n526) );
  NAND2_X2 U903 ( .A1(regBoiz_regfile_26__20_), .A2(n6742), .ZN(n527) );
  NAND2_X2 U905 ( .A1(regBoiz_regfile_26__1_), .A2(n6742), .ZN(n528) );
  NAND2_X2 U907 ( .A1(regBoiz_regfile_26__19_), .A2(n6742), .ZN(n529) );
  NAND2_X2 U909 ( .A1(regBoiz_regfile_26__18_), .A2(n6742), .ZN(n530) );
  NAND2_X2 U911 ( .A1(regBoiz_regfile_26__17_), .A2(n6742), .ZN(n531) );
  NAND2_X2 U913 ( .A1(regBoiz_regfile_26__16_), .A2(n507), .ZN(n532) );
  NAND2_X2 U915 ( .A1(regBoiz_regfile_26__15_), .A2(n6741), .ZN(n533) );
  NAND2_X2 U917 ( .A1(regBoiz_regfile_26__14_), .A2(n6742), .ZN(n534) );
  NAND2_X2 U919 ( .A1(regBoiz_regfile_26__13_), .A2(n507), .ZN(n535) );
  NAND2_X2 U921 ( .A1(regBoiz_regfile_26__12_), .A2(n6742), .ZN(n536) );
  NAND2_X2 U923 ( .A1(regBoiz_regfile_26__11_), .A2(n6742), .ZN(n537) );
  NAND2_X2 U927 ( .A1(regBoiz_regfile_26__0_), .A2(n6742), .ZN(n539) );
  NAND2_X2 U928 ( .A1(n506), .A2(n203), .ZN(n507) );
  NAND2_X2 U932 ( .A1(regBoiz_regfile_25__8_), .A2(n6736), .ZN(n542) );
  NAND2_X2 U934 ( .A1(regBoiz_regfile_25__7_), .A2(n6737), .ZN(n543) );
  NAND2_X2 U936 ( .A1(regBoiz_regfile_25__6_), .A2(n6736), .ZN(n544) );
  NAND2_X2 U938 ( .A1(regBoiz_regfile_25__5_), .A2(n6737), .ZN(n545) );
  NAND2_X2 U942 ( .A1(regBoiz_regfile_25__3_), .A2(n6736), .ZN(n547) );
  NAND2_X2 U944 ( .A1(regBoiz_regfile_25__31_), .A2(n6737), .ZN(n548) );
  NAND2_X2 U946 ( .A1(regBoiz_regfile_25__30_), .A2(n6738), .ZN(n549) );
  NAND2_X2 U948 ( .A1(regBoiz_regfile_25__2_), .A2(n6738), .ZN(n550) );
  NAND2_X2 U950 ( .A1(regBoiz_regfile_25__29_), .A2(n6738), .ZN(n551) );
  NAND2_X2 U952 ( .A1(regBoiz_regfile_25__28_), .A2(n6738), .ZN(n552) );
  NAND2_X2 U954 ( .A1(regBoiz_regfile_25__27_), .A2(n6738), .ZN(n553) );
  NAND2_X2 U956 ( .A1(regBoiz_regfile_25__26_), .A2(n6738), .ZN(n554) );
  NAND2_X2 U958 ( .A1(regBoiz_regfile_25__25_), .A2(n6738), .ZN(n555) );
  NAND2_X2 U960 ( .A1(regBoiz_regfile_25__24_), .A2(n6738), .ZN(n556) );
  NAND2_X2 U962 ( .A1(regBoiz_regfile_25__23_), .A2(n6738), .ZN(n557) );
  NAND2_X2 U964 ( .A1(regBoiz_regfile_25__22_), .A2(n6738), .ZN(n558) );
  NAND2_X2 U966 ( .A1(regBoiz_regfile_25__21_), .A2(n6738), .ZN(n559) );
  NAND2_X2 U968 ( .A1(regBoiz_regfile_25__20_), .A2(n6738), .ZN(n560) );
  NAND2_X2 U970 ( .A1(regBoiz_regfile_25__1_), .A2(n6738), .ZN(n561) );
  NAND2_X2 U972 ( .A1(regBoiz_regfile_25__19_), .A2(n6738), .ZN(n562) );
  NAND2_X2 U974 ( .A1(regBoiz_regfile_25__18_), .A2(n6738), .ZN(n563) );
  NAND2_X2 U976 ( .A1(regBoiz_regfile_25__17_), .A2(n6738), .ZN(n564) );
  NAND2_X2 U978 ( .A1(regBoiz_regfile_25__16_), .A2(n540), .ZN(n565) );
  NAND2_X2 U980 ( .A1(regBoiz_regfile_25__15_), .A2(n6737), .ZN(n566) );
  NAND2_X2 U982 ( .A1(regBoiz_regfile_25__14_), .A2(n6738), .ZN(n567) );
  NAND2_X2 U984 ( .A1(regBoiz_regfile_25__13_), .A2(n6736), .ZN(n568) );
  NAND2_X2 U986 ( .A1(regBoiz_regfile_25__12_), .A2(n6738), .ZN(n569) );
  NAND2_X2 U988 ( .A1(regBoiz_regfile_25__11_), .A2(n6738), .ZN(n570) );
  NAND2_X2 U992 ( .A1(regBoiz_regfile_25__0_), .A2(n6738), .ZN(n572) );
  NAND2_X2 U993 ( .A1(n506), .A2(n99), .ZN(n540) );
  NAND2_X2 U995 ( .A1(regBoiz_regfile_24__9_), .A2(n6734), .ZN(n574) );
  NAND2_X2 U997 ( .A1(regBoiz_regfile_24__8_), .A2(n6733), .ZN(n575) );
  NAND2_X2 U999 ( .A1(regBoiz_regfile_24__7_), .A2(n6732), .ZN(n576) );
  NAND2_X2 U1001 ( .A1(regBoiz_regfile_24__6_), .A2(n6733), .ZN(n577) );
  NAND2_X2 U1003 ( .A1(regBoiz_regfile_24__5_), .A2(n6732), .ZN(n578) );
  NAND2_X2 U1005 ( .A1(regBoiz_regfile_24__4_), .A2(n6733), .ZN(n579) );
  NAND2_X2 U1007 ( .A1(regBoiz_regfile_24__3_), .A2(n6732), .ZN(n580) );
  NAND2_X2 U1009 ( .A1(regBoiz_regfile_24__31_), .A2(n6734), .ZN(n581) );
  NAND2_X2 U1011 ( .A1(regBoiz_regfile_24__30_), .A2(n6732), .ZN(n582) );
  NAND2_X2 U1013 ( .A1(regBoiz_regfile_24__2_), .A2(n6733), .ZN(n583) );
  NAND2_X2 U1015 ( .A1(regBoiz_regfile_24__29_), .A2(n6734), .ZN(n584) );
  NAND2_X2 U1019 ( .A1(regBoiz_regfile_24__27_), .A2(n6734), .ZN(n586) );
  NAND2_X2 U1021 ( .A1(regBoiz_regfile_24__26_), .A2(n573), .ZN(n587) );
  NAND2_X2 U1023 ( .A1(regBoiz_regfile_24__25_), .A2(n573), .ZN(n588) );
  NAND2_X2 U1025 ( .A1(regBoiz_regfile_24__24_), .A2(n573), .ZN(n589) );
  NAND2_X2 U1027 ( .A1(regBoiz_regfile_24__23_), .A2(n573), .ZN(n590) );
  NAND2_X2 U1029 ( .A1(regBoiz_regfile_24__22_), .A2(n573), .ZN(n591) );
  NAND2_X2 U1031 ( .A1(regBoiz_regfile_24__21_), .A2(n6734), .ZN(n592) );
  NAND2_X2 U1033 ( .A1(regBoiz_regfile_24__20_), .A2(n573), .ZN(n593) );
  NAND2_X2 U1035 ( .A1(regBoiz_regfile_24__1_), .A2(n573), .ZN(n594) );
  NAND2_X2 U1037 ( .A1(regBoiz_regfile_24__19_), .A2(n573), .ZN(n595) );
  NAND2_X2 U1039 ( .A1(regBoiz_regfile_24__18_), .A2(n6734), .ZN(n596) );
  NAND2_X2 U1041 ( .A1(regBoiz_regfile_24__17_), .A2(n573), .ZN(n597) );
  NAND2_X2 U1043 ( .A1(regBoiz_regfile_24__16_), .A2(n6734), .ZN(n598) );
  NAND2_X2 U1045 ( .A1(regBoiz_regfile_24__15_), .A2(n6734), .ZN(n599) );
  NAND2_X2 U1047 ( .A1(regBoiz_regfile_24__14_), .A2(n573), .ZN(n600) );
  NAND2_X2 U1049 ( .A1(regBoiz_regfile_24__13_), .A2(n6734), .ZN(n601) );
  NAND2_X2 U1051 ( .A1(regBoiz_regfile_24__12_), .A2(n6734), .ZN(n602) );
  NAND2_X2 U1053 ( .A1(regBoiz_regfile_24__11_), .A2(n573), .ZN(n603) );
  NAND2_X2 U1055 ( .A1(regBoiz_regfile_24__10_), .A2(n6734), .ZN(n604) );
  NAND2_X2 U1057 ( .A1(regBoiz_regfile_24__0_), .A2(n573), .ZN(n605) );
  NAND2_X2 U1058 ( .A1(n506), .A2(n134), .ZN(n573) );
  AND2_X2 U1059 ( .A1(n472), .A2(n5482), .ZN(n506) );
  AND2_X2 U1060 ( .A1(n607), .A2(wbRwh[3]), .ZN(n472) );
  NAND2_X2 U1062 ( .A1(regBoiz_regfile_23__9_), .A2(n6730), .ZN(n609) );
  NAND2_X2 U1064 ( .A1(regBoiz_regfile_23__8_), .A2(n6728), .ZN(n610) );
  NAND2_X2 U1066 ( .A1(regBoiz_regfile_23__7_), .A2(n6729), .ZN(n611) );
  NAND2_X2 U1070 ( .A1(regBoiz_regfile_23__5_), .A2(n6729), .ZN(n613) );
  NAND2_X2 U1072 ( .A1(regBoiz_regfile_23__4_), .A2(n6728), .ZN(n614) );
  NAND2_X2 U1074 ( .A1(regBoiz_regfile_23__3_), .A2(n6729), .ZN(n615) );
  NAND2_X2 U1076 ( .A1(regBoiz_regfile_23__31_), .A2(n6728), .ZN(n616) );
  NAND2_X2 U1078 ( .A1(regBoiz_regfile_23__30_), .A2(n6730), .ZN(n617) );
  NAND2_X2 U1080 ( .A1(regBoiz_regfile_23__2_), .A2(n6730), .ZN(n618) );
  NAND2_X2 U1082 ( .A1(regBoiz_regfile_23__29_), .A2(n6730), .ZN(n619) );
  NAND2_X2 U1084 ( .A1(regBoiz_regfile_23__28_), .A2(n6730), .ZN(n620) );
  NAND2_X2 U1086 ( .A1(regBoiz_regfile_23__27_), .A2(n6730), .ZN(n621) );
  NAND2_X2 U1088 ( .A1(regBoiz_regfile_23__26_), .A2(n6730), .ZN(n622) );
  NAND2_X2 U1090 ( .A1(regBoiz_regfile_23__25_), .A2(n6730), .ZN(n623) );
  NAND2_X2 U1092 ( .A1(regBoiz_regfile_23__24_), .A2(n6730), .ZN(n624) );
  NAND2_X2 U1096 ( .A1(regBoiz_regfile_23__22_), .A2(n6730), .ZN(n626) );
  NAND2_X2 U1098 ( .A1(regBoiz_regfile_23__21_), .A2(n6730), .ZN(n627) );
  NAND2_X2 U1100 ( .A1(regBoiz_regfile_23__20_), .A2(n6730), .ZN(n628) );
  NAND2_X2 U1104 ( .A1(regBoiz_regfile_23__19_), .A2(n6730), .ZN(n630) );
  NAND2_X2 U1106 ( .A1(regBoiz_regfile_23__18_), .A2(n6730), .ZN(n631) );
  NAND2_X2 U1108 ( .A1(regBoiz_regfile_23__17_), .A2(n6730), .ZN(n632) );
  NAND2_X2 U1110 ( .A1(regBoiz_regfile_23__16_), .A2(n6730), .ZN(n633) );
  NAND2_X2 U1112 ( .A1(regBoiz_regfile_23__15_), .A2(n6730), .ZN(n634) );
  NAND2_X2 U1114 ( .A1(regBoiz_regfile_23__14_), .A2(n6730), .ZN(n635) );
  NAND2_X2 U1116 ( .A1(regBoiz_regfile_23__13_), .A2(n6730), .ZN(n636) );
  NAND2_X2 U1118 ( .A1(regBoiz_regfile_23__12_), .A2(n6730), .ZN(n637) );
  NAND2_X2 U1120 ( .A1(regBoiz_regfile_23__11_), .A2(n6730), .ZN(n638) );
  NAND2_X2 U1124 ( .A1(regBoiz_regfile_23__0_), .A2(n6730), .ZN(n640) );
  NAND2_X2 U1127 ( .A1(regBoiz_regfile_22__9_), .A2(n6727), .ZN(n643) );
  NAND2_X2 U1129 ( .A1(regBoiz_regfile_22__8_), .A2(n6726), .ZN(n644) );
  NAND2_X2 U1131 ( .A1(regBoiz_regfile_22__7_), .A2(n6725), .ZN(n645) );
  NAND2_X2 U1133 ( .A1(regBoiz_regfile_22__6_), .A2(n6726), .ZN(n646) );
  NAND2_X2 U1135 ( .A1(regBoiz_regfile_22__5_), .A2(n6725), .ZN(n647) );
  NAND2_X2 U1137 ( .A1(regBoiz_regfile_22__4_), .A2(n6725), .ZN(n648) );
  NAND2_X2 U1139 ( .A1(regBoiz_regfile_22__3_), .A2(n6726), .ZN(n649) );
  NAND2_X2 U1141 ( .A1(regBoiz_regfile_22__31_), .A2(n6725), .ZN(n650) );
  NAND2_X2 U1143 ( .A1(regBoiz_regfile_22__30_), .A2(n6727), .ZN(n651) );
  NAND2_X2 U1145 ( .A1(regBoiz_regfile_22__2_), .A2(n6727), .ZN(n652) );
  NAND2_X2 U1147 ( .A1(regBoiz_regfile_22__29_), .A2(n6727), .ZN(n653) );
  NAND2_X2 U1151 ( .A1(regBoiz_regfile_22__27_), .A2(n6727), .ZN(n655) );
  NAND2_X2 U1153 ( .A1(regBoiz_regfile_22__26_), .A2(n6727), .ZN(n656) );
  NAND2_X2 U1155 ( .A1(regBoiz_regfile_22__25_), .A2(n6727), .ZN(n657) );
  NAND2_X2 U1157 ( .A1(regBoiz_regfile_22__24_), .A2(n6727), .ZN(n658) );
  NAND2_X2 U1159 ( .A1(regBoiz_regfile_22__23_), .A2(n6727), .ZN(n659) );
  NAND2_X2 U1161 ( .A1(regBoiz_regfile_22__22_), .A2(n6727), .ZN(n660) );
  NAND2_X2 U1163 ( .A1(regBoiz_regfile_22__21_), .A2(n6727), .ZN(n661) );
  NAND2_X2 U1165 ( .A1(regBoiz_regfile_22__20_), .A2(n6727), .ZN(n662) );
  NAND2_X2 U1167 ( .A1(regBoiz_regfile_22__1_), .A2(n6727), .ZN(n663) );
  NAND2_X2 U1169 ( .A1(regBoiz_regfile_22__19_), .A2(n6727), .ZN(n664) );
  NAND2_X2 U1171 ( .A1(regBoiz_regfile_22__18_), .A2(n6727), .ZN(n665) );
  NAND2_X2 U1173 ( .A1(regBoiz_regfile_22__17_), .A2(n6727), .ZN(n666) );
  NAND2_X2 U1175 ( .A1(regBoiz_regfile_22__16_), .A2(n6727), .ZN(n667) );
  NAND2_X2 U1177 ( .A1(regBoiz_regfile_22__15_), .A2(n6727), .ZN(n668) );
  NAND2_X2 U1179 ( .A1(regBoiz_regfile_22__14_), .A2(n6727), .ZN(n669) );
  NAND2_X2 U1181 ( .A1(regBoiz_regfile_22__13_), .A2(n6727), .ZN(n670) );
  NAND2_X2 U1183 ( .A1(regBoiz_regfile_22__12_), .A2(n6727), .ZN(n671) );
  NAND2_X2 U1185 ( .A1(regBoiz_regfile_22__11_), .A2(n6727), .ZN(n672) );
  NAND2_X2 U1189 ( .A1(regBoiz_regfile_22__0_), .A2(n6727), .ZN(n674) );
  NAND2_X2 U1194 ( .A1(regBoiz_regfile_21__8_), .A2(n6723), .ZN(n677) );
  NAND2_X2 U1196 ( .A1(regBoiz_regfile_21__7_), .A2(n6722), .ZN(n678) );
  NAND2_X2 U1198 ( .A1(regBoiz_regfile_21__6_), .A2(n6723), .ZN(n679) );
  NAND2_X2 U1200 ( .A1(regBoiz_regfile_21__5_), .A2(n6722), .ZN(n680) );
  NAND2_X2 U1202 ( .A1(regBoiz_regfile_21__4_), .A2(n6722), .ZN(n681) );
  NAND2_X2 U1204 ( .A1(regBoiz_regfile_21__3_), .A2(n6723), .ZN(n682) );
  NAND2_X2 U1206 ( .A1(regBoiz_regfile_21__31_), .A2(n6724), .ZN(n683) );
  NAND2_X2 U1208 ( .A1(regBoiz_regfile_21__30_), .A2(n6724), .ZN(n684) );
  NAND2_X2 U1210 ( .A1(regBoiz_regfile_21__2_), .A2(n6724), .ZN(n685) );
  NAND2_X2 U1212 ( .A1(regBoiz_regfile_21__29_), .A2(n6724), .ZN(n686) );
  NAND2_X2 U1214 ( .A1(regBoiz_regfile_21__28_), .A2(n6724), .ZN(n687) );
  NAND2_X2 U1216 ( .A1(regBoiz_regfile_21__27_), .A2(n6724), .ZN(n688) );
  NAND2_X2 U1218 ( .A1(regBoiz_regfile_21__26_), .A2(n6724), .ZN(n689) );
  NAND2_X2 U1220 ( .A1(regBoiz_regfile_21__25_), .A2(n6724), .ZN(n690) );
  NAND2_X2 U1222 ( .A1(regBoiz_regfile_21__24_), .A2(n6724), .ZN(n691) );
  NAND2_X2 U1224 ( .A1(regBoiz_regfile_21__23_), .A2(n6724), .ZN(n692) );
  NAND2_X2 U1226 ( .A1(regBoiz_regfile_21__22_), .A2(n6724), .ZN(n693) );
  NAND2_X2 U1228 ( .A1(regBoiz_regfile_21__21_), .A2(n6724), .ZN(n694) );
  NAND2_X2 U1230 ( .A1(regBoiz_regfile_21__20_), .A2(n6724), .ZN(n695) );
  NAND2_X2 U1232 ( .A1(regBoiz_regfile_21__1_), .A2(n6724), .ZN(n696) );
  NAND2_X2 U1234 ( .A1(regBoiz_regfile_21__19_), .A2(n6724), .ZN(n697) );
  NAND2_X2 U1236 ( .A1(regBoiz_regfile_21__18_), .A2(n6724), .ZN(n698) );
  NAND2_X2 U1238 ( .A1(regBoiz_regfile_21__17_), .A2(n6724), .ZN(n699) );
  NAND2_X2 U1240 ( .A1(regBoiz_regfile_21__16_), .A2(n6723), .ZN(n700) );
  NAND2_X2 U1242 ( .A1(regBoiz_regfile_21__15_), .A2(n6724), .ZN(n701) );
  NAND2_X2 U1244 ( .A1(regBoiz_regfile_21__14_), .A2(n6724), .ZN(n702) );
  NAND2_X2 U1246 ( .A1(regBoiz_regfile_21__13_), .A2(n6722), .ZN(n703) );
  NAND2_X2 U1248 ( .A1(regBoiz_regfile_21__12_), .A2(n6724), .ZN(n704) );
  NAND2_X2 U1250 ( .A1(regBoiz_regfile_21__11_), .A2(n6724), .ZN(n705) );
  NAND2_X2 U1252 ( .A1(regBoiz_regfile_21__10_), .A2(n6724), .ZN(n706) );
  NAND2_X2 U1254 ( .A1(regBoiz_regfile_21__0_), .A2(n6724), .ZN(n707) );
  NAND2_X2 U1255 ( .A1(n641), .A2(n99), .ZN(n675) );
  NAND2_X2 U1257 ( .A1(regBoiz_regfile_20__9_), .A2(n6719), .ZN(n709) );
  NAND2_X2 U1259 ( .A1(regBoiz_regfile_20__8_), .A2(n6718), .ZN(n710) );
  NAND2_X2 U1261 ( .A1(regBoiz_regfile_20__7_), .A2(n6717), .ZN(n711) );
  NAND2_X2 U1263 ( .A1(regBoiz_regfile_20__6_), .A2(n6718), .ZN(n712) );
  NAND2_X2 U1265 ( .A1(regBoiz_regfile_20__5_), .A2(n6717), .ZN(n713) );
  NAND2_X2 U1267 ( .A1(regBoiz_regfile_20__4_), .A2(n6717), .ZN(n714) );
  NAND2_X2 U1269 ( .A1(regBoiz_regfile_20__3_), .A2(n6718), .ZN(n715) );
  NAND2_X2 U1271 ( .A1(regBoiz_regfile_20__31_), .A2(n6719), .ZN(n716) );
  NAND2_X2 U1273 ( .A1(regBoiz_regfile_20__30_), .A2(n6719), .ZN(n717) );
  NAND2_X2 U1275 ( .A1(regBoiz_regfile_20__2_), .A2(n6719), .ZN(n718) );
  NAND2_X2 U1277 ( .A1(regBoiz_regfile_20__29_), .A2(n6719), .ZN(n719) );
  NAND2_X2 U1279 ( .A1(regBoiz_regfile_20__28_), .A2(n6719), .ZN(n720) );
  NAND2_X2 U1281 ( .A1(regBoiz_regfile_20__27_), .A2(n6719), .ZN(n721) );
  NAND2_X2 U1283 ( .A1(regBoiz_regfile_20__26_), .A2(n6719), .ZN(n722) );
  NAND2_X2 U1285 ( .A1(regBoiz_regfile_20__25_), .A2(n6719), .ZN(n723) );
  NAND2_X2 U1287 ( .A1(regBoiz_regfile_20__24_), .A2(n6719), .ZN(n724) );
  NAND2_X2 U1289 ( .A1(regBoiz_regfile_20__23_), .A2(n6719), .ZN(n725) );
  NAND2_X2 U1291 ( .A1(regBoiz_regfile_20__22_), .A2(n6719), .ZN(n726) );
  NAND2_X2 U1293 ( .A1(regBoiz_regfile_20__21_), .A2(n6719), .ZN(n727) );
  NAND2_X2 U1295 ( .A1(regBoiz_regfile_20__20_), .A2(n6719), .ZN(n728) );
  NAND2_X2 U1297 ( .A1(regBoiz_regfile_20__1_), .A2(n6719), .ZN(n729) );
  NAND2_X2 U1299 ( .A1(regBoiz_regfile_20__19_), .A2(n6719), .ZN(n730) );
  NAND2_X2 U1301 ( .A1(regBoiz_regfile_20__18_), .A2(n6719), .ZN(n731) );
  NAND2_X2 U1303 ( .A1(regBoiz_regfile_20__17_), .A2(n6719), .ZN(n732) );
  NAND2_X2 U1305 ( .A1(regBoiz_regfile_20__16_), .A2(n708), .ZN(n733) );
  NAND2_X2 U1307 ( .A1(regBoiz_regfile_20__15_), .A2(n6718), .ZN(n734) );
  NAND2_X2 U1309 ( .A1(regBoiz_regfile_20__14_), .A2(n6719), .ZN(n735) );
  NAND2_X2 U1311 ( .A1(regBoiz_regfile_20__13_), .A2(n6717), .ZN(n736) );
  NAND2_X2 U1313 ( .A1(regBoiz_regfile_20__12_), .A2(n6719), .ZN(n737) );
  NAND2_X2 U1315 ( .A1(regBoiz_regfile_20__11_), .A2(n6719), .ZN(n738) );
  NAND2_X2 U1317 ( .A1(regBoiz_regfile_20__10_), .A2(n6719), .ZN(n739) );
  NAND2_X2 U1319 ( .A1(regBoiz_regfile_20__0_), .A2(n6719), .ZN(n740) );
  NAND2_X2 U1320 ( .A1(n641), .A2(n134), .ZN(n708) );
  AND2_X2 U1321 ( .A1(n607), .A2(n270), .ZN(n641) );
  NAND2_X2 U1324 ( .A1(regBoiz_regfile_1__9_), .A2(n6715), .ZN(n742) );
  NAND2_X2 U1326 ( .A1(regBoiz_regfile_1__8_), .A2(n6713), .ZN(n743) );
  NAND2_X2 U1328 ( .A1(regBoiz_regfile_1__7_), .A2(n6714), .ZN(n744) );
  NAND2_X2 U1330 ( .A1(regBoiz_regfile_1__6_), .A2(n6713), .ZN(n745) );
  NAND2_X2 U1332 ( .A1(regBoiz_regfile_1__5_), .A2(n6714), .ZN(n746) );
  NAND2_X2 U1334 ( .A1(regBoiz_regfile_1__4_), .A2(n6713), .ZN(n747) );
  NAND2_X2 U1336 ( .A1(regBoiz_regfile_1__3_), .A2(n6714), .ZN(n748) );
  NAND2_X2 U1338 ( .A1(regBoiz_regfile_1__31_), .A2(n6715), .ZN(n749) );
  NAND2_X2 U1340 ( .A1(regBoiz_regfile_1__30_), .A2(n6715), .ZN(n750) );
  NAND2_X2 U1342 ( .A1(regBoiz_regfile_1__2_), .A2(n6715), .ZN(n751) );
  NAND2_X2 U1344 ( .A1(regBoiz_regfile_1__29_), .A2(n6715), .ZN(n752) );
  NAND2_X2 U1346 ( .A1(regBoiz_regfile_1__28_), .A2(n6715), .ZN(n753) );
  NAND2_X2 U1348 ( .A1(regBoiz_regfile_1__27_), .A2(n6715), .ZN(n754) );
  NAND2_X2 U1350 ( .A1(regBoiz_regfile_1__26_), .A2(n6715), .ZN(n755) );
  NAND2_X2 U1352 ( .A1(regBoiz_regfile_1__25_), .A2(n6715), .ZN(n756) );
  NAND2_X2 U1354 ( .A1(regBoiz_regfile_1__24_), .A2(n6715), .ZN(n757) );
  NAND2_X2 U1356 ( .A1(regBoiz_regfile_1__23_), .A2(n6715), .ZN(n758) );
  NAND2_X2 U1358 ( .A1(regBoiz_regfile_1__22_), .A2(n6715), .ZN(n759) );
  NAND2_X2 U1360 ( .A1(regBoiz_regfile_1__21_), .A2(n6715), .ZN(n760) );
  NAND2_X2 U1362 ( .A1(regBoiz_regfile_1__20_), .A2(n6715), .ZN(n761) );
  NAND2_X2 U1364 ( .A1(regBoiz_regfile_1__1_), .A2(n6715), .ZN(n762) );
  NAND2_X2 U1366 ( .A1(regBoiz_regfile_1__19_), .A2(n6715), .ZN(n763) );
  NAND2_X2 U1368 ( .A1(regBoiz_regfile_1__18_), .A2(n6715), .ZN(n764) );
  NAND2_X2 U1370 ( .A1(regBoiz_regfile_1__17_), .A2(n6715), .ZN(n765) );
  NAND2_X2 U1372 ( .A1(regBoiz_regfile_1__16_), .A2(n6715), .ZN(n766) );
  NAND2_X2 U1374 ( .A1(regBoiz_regfile_1__15_), .A2(n6714), .ZN(n767) );
  NAND2_X2 U1376 ( .A1(regBoiz_regfile_1__14_), .A2(n6715), .ZN(n768) );
  NAND2_X2 U1378 ( .A1(regBoiz_regfile_1__13_), .A2(n6713), .ZN(n769) );
  NAND2_X2 U1380 ( .A1(regBoiz_regfile_1__12_), .A2(n6715), .ZN(n770) );
  NAND2_X2 U1382 ( .A1(regBoiz_regfile_1__11_), .A2(n6715), .ZN(n771) );
  NAND2_X2 U1384 ( .A1(regBoiz_regfile_1__10_), .A2(n6715), .ZN(n772) );
  NAND2_X2 U1386 ( .A1(regBoiz_regfile_1__0_), .A2(n6715), .ZN(n773) );
  NAND2_X2 U1387 ( .A1(n305), .A2(n99), .ZN(n741) );
  NAND2_X2 U1389 ( .A1(regBoiz_regfile_19__9_), .A2(n6712), .ZN(n775) );
  NAND2_X2 U1391 ( .A1(regBoiz_regfile_19__8_), .A2(n6710), .ZN(n776) );
  NAND2_X2 U1393 ( .A1(regBoiz_regfile_19__7_), .A2(n6711), .ZN(n777) );
  NAND2_X2 U1395 ( .A1(regBoiz_regfile_19__6_), .A2(n6710), .ZN(n778) );
  NAND2_X2 U1397 ( .A1(regBoiz_regfile_19__5_), .A2(n6711), .ZN(n779) );
  NAND2_X2 U1399 ( .A1(regBoiz_regfile_19__4_), .A2(n6711), .ZN(n780) );
  NAND2_X2 U1401 ( .A1(regBoiz_regfile_19__3_), .A2(n6710), .ZN(n781) );
  NAND2_X2 U1403 ( .A1(regBoiz_regfile_19__31_), .A2(n6711), .ZN(n782) );
  NAND2_X2 U1405 ( .A1(regBoiz_regfile_19__30_), .A2(n6712), .ZN(n783) );
  NAND2_X2 U1407 ( .A1(regBoiz_regfile_19__2_), .A2(n6712), .ZN(n784) );
  NAND2_X2 U1409 ( .A1(regBoiz_regfile_19__29_), .A2(n6712), .ZN(n785) );
  NAND2_X2 U1413 ( .A1(regBoiz_regfile_19__27_), .A2(n6712), .ZN(n787) );
  NAND2_X2 U1415 ( .A1(regBoiz_regfile_19__26_), .A2(n6712), .ZN(n788) );
  NAND2_X2 U1417 ( .A1(regBoiz_regfile_19__25_), .A2(n6712), .ZN(n789) );
  NAND2_X2 U1419 ( .A1(regBoiz_regfile_19__24_), .A2(n6712), .ZN(n790) );
  NAND2_X2 U1421 ( .A1(regBoiz_regfile_19__23_), .A2(n6712), .ZN(n791) );
  NAND2_X2 U1423 ( .A1(regBoiz_regfile_19__22_), .A2(n6712), .ZN(n792) );
  NAND2_X2 U1425 ( .A1(regBoiz_regfile_19__21_), .A2(n6712), .ZN(n793) );
  NAND2_X2 U1427 ( .A1(regBoiz_regfile_19__20_), .A2(n6712), .ZN(n794) );
  NAND2_X2 U1429 ( .A1(regBoiz_regfile_19__1_), .A2(n6712), .ZN(n795) );
  NAND2_X2 U1431 ( .A1(regBoiz_regfile_19__19_), .A2(n6712), .ZN(n796) );
  NAND2_X2 U1433 ( .A1(regBoiz_regfile_19__18_), .A2(n6712), .ZN(n797) );
  NAND2_X2 U1435 ( .A1(regBoiz_regfile_19__17_), .A2(n6712), .ZN(n798) );
  NAND2_X2 U1437 ( .A1(regBoiz_regfile_19__16_), .A2(n6712), .ZN(n799) );
  NAND2_X2 U1439 ( .A1(regBoiz_regfile_19__15_), .A2(n6712), .ZN(n800) );
  NAND2_X2 U1441 ( .A1(regBoiz_regfile_19__14_), .A2(n6712), .ZN(n801) );
  NAND2_X2 U1443 ( .A1(regBoiz_regfile_19__13_), .A2(n6712), .ZN(n802) );
  NAND2_X2 U1445 ( .A1(regBoiz_regfile_19__12_), .A2(n6712), .ZN(n803) );
  NAND2_X2 U1447 ( .A1(regBoiz_regfile_19__11_), .A2(n6712), .ZN(n804) );
  NAND2_X2 U1451 ( .A1(regBoiz_regfile_19__0_), .A2(n6712), .ZN(n806) );
  NAND2_X2 U1454 ( .A1(regBoiz_regfile_18__9_), .A2(n6709), .ZN(n809) );
  NAND2_X2 U1456 ( .A1(regBoiz_regfile_18__8_), .A2(n6708), .ZN(n810) );
  NAND2_X2 U1458 ( .A1(regBoiz_regfile_18__7_), .A2(n6707), .ZN(n811) );
  NAND2_X2 U1460 ( .A1(regBoiz_regfile_18__6_), .A2(n6708), .ZN(n812) );
  NAND2_X2 U1462 ( .A1(regBoiz_regfile_18__5_), .A2(n6707), .ZN(n813) );
  NAND2_X2 U1464 ( .A1(regBoiz_regfile_18__4_), .A2(n6708), .ZN(n814) );
  NAND2_X2 U1466 ( .A1(regBoiz_regfile_18__3_), .A2(n6707), .ZN(n815) );
  NAND2_X2 U1468 ( .A1(regBoiz_regfile_18__31_), .A2(n6708), .ZN(n816) );
  NAND2_X2 U1470 ( .A1(regBoiz_regfile_18__30_), .A2(n6709), .ZN(n817) );
  NAND2_X2 U1472 ( .A1(regBoiz_regfile_18__2_), .A2(n6709), .ZN(n818) );
  NAND2_X2 U1474 ( .A1(regBoiz_regfile_18__29_), .A2(n6709), .ZN(n819) );
  NAND2_X2 U1478 ( .A1(regBoiz_regfile_18__27_), .A2(n6709), .ZN(n821) );
  NAND2_X2 U1480 ( .A1(regBoiz_regfile_18__26_), .A2(n6709), .ZN(n822) );
  NAND2_X2 U1482 ( .A1(regBoiz_regfile_18__25_), .A2(n6709), .ZN(n823) );
  NAND2_X2 U1484 ( .A1(regBoiz_regfile_18__24_), .A2(n6709), .ZN(n824) );
  NAND2_X2 U1486 ( .A1(regBoiz_regfile_18__23_), .A2(n6709), .ZN(n825) );
  NAND2_X2 U1488 ( .A1(regBoiz_regfile_18__22_), .A2(n6709), .ZN(n826) );
  NAND2_X2 U1490 ( .A1(regBoiz_regfile_18__21_), .A2(n6709), .ZN(n827) );
  NAND2_X2 U1492 ( .A1(regBoiz_regfile_18__20_), .A2(n6709), .ZN(n828) );
  NAND2_X2 U1494 ( .A1(regBoiz_regfile_18__1_), .A2(n6709), .ZN(n829) );
  NAND2_X2 U1496 ( .A1(regBoiz_regfile_18__19_), .A2(n6709), .ZN(n830) );
  NAND2_X2 U1498 ( .A1(regBoiz_regfile_18__18_), .A2(n6709), .ZN(n831) );
  NAND2_X2 U1500 ( .A1(regBoiz_regfile_18__17_), .A2(n6709), .ZN(n832) );
  NAND2_X2 U1502 ( .A1(regBoiz_regfile_18__16_), .A2(n6709), .ZN(n833) );
  NAND2_X2 U1504 ( .A1(regBoiz_regfile_18__15_), .A2(n6709), .ZN(n834) );
  NAND2_X2 U1506 ( .A1(regBoiz_regfile_18__14_), .A2(n6709), .ZN(n835) );
  NAND2_X2 U1508 ( .A1(regBoiz_regfile_18__13_), .A2(n6709), .ZN(n836) );
  NAND2_X2 U1510 ( .A1(regBoiz_regfile_18__12_), .A2(n6709), .ZN(n837) );
  NAND2_X2 U1512 ( .A1(regBoiz_regfile_18__11_), .A2(n6709), .ZN(n838) );
  NAND2_X2 U1514 ( .A1(regBoiz_regfile_18__10_), .A2(n6709), .ZN(n839) );
  NAND2_X2 U1516 ( .A1(regBoiz_regfile_18__0_), .A2(n6709), .ZN(n840) );
  NAND2_X2 U1519 ( .A1(regBoiz_regfile_17__9_), .A2(n6706), .ZN(n842) );
  NAND2_X2 U1521 ( .A1(regBoiz_regfile_17__8_), .A2(n6705), .ZN(n843) );
  NAND2_X2 U1523 ( .A1(regBoiz_regfile_17__7_), .A2(n6705), .ZN(n844) );
  NAND2_X2 U1525 ( .A1(regBoiz_regfile_17__6_), .A2(n6705), .ZN(n845) );
  NAND2_X2 U1527 ( .A1(regBoiz_regfile_17__5_), .A2(n6705), .ZN(n846) );
  NAND2_X2 U1531 ( .A1(regBoiz_regfile_17__3_), .A2(n6706), .ZN(n848) );
  NAND2_X2 U1533 ( .A1(regBoiz_regfile_17__31_), .A2(n6705), .ZN(n849) );
  NAND2_X2 U1535 ( .A1(regBoiz_regfile_17__30_), .A2(n6704), .ZN(n850) );
  NAND2_X2 U1537 ( .A1(regBoiz_regfile_17__2_), .A2(n6706), .ZN(n851) );
  NAND2_X2 U1539 ( .A1(regBoiz_regfile_17__29_), .A2(n6706), .ZN(n852) );
  NAND2_X2 U1543 ( .A1(regBoiz_regfile_17__27_), .A2(n6704), .ZN(n854) );
  NAND2_X2 U1545 ( .A1(regBoiz_regfile_17__26_), .A2(n6706), .ZN(n855) );
  NAND2_X2 U1547 ( .A1(regBoiz_regfile_17__25_), .A2(n6704), .ZN(n856) );
  NAND2_X2 U1549 ( .A1(regBoiz_regfile_17__24_), .A2(n6706), .ZN(n857) );
  NAND2_X2 U1551 ( .A1(regBoiz_regfile_17__23_), .A2(n6704), .ZN(n858) );
  NAND2_X2 U1553 ( .A1(regBoiz_regfile_17__22_), .A2(n841), .ZN(n859) );
  NAND2_X2 U1555 ( .A1(regBoiz_regfile_17__21_), .A2(n6706), .ZN(n860) );
  NAND2_X2 U1557 ( .A1(regBoiz_regfile_17__20_), .A2(n841), .ZN(n861) );
  NAND2_X2 U1559 ( .A1(regBoiz_regfile_17__1_), .A2(n841), .ZN(n862) );
  NAND2_X2 U1561 ( .A1(regBoiz_regfile_17__19_), .A2(n841), .ZN(n863) );
  NAND2_X2 U1563 ( .A1(regBoiz_regfile_17__18_), .A2(n6706), .ZN(n864) );
  NAND2_X2 U1565 ( .A1(regBoiz_regfile_17__17_), .A2(n841), .ZN(n865) );
  NAND2_X2 U1567 ( .A1(regBoiz_regfile_17__16_), .A2(n6706), .ZN(n866) );
  NAND2_X2 U1569 ( .A1(regBoiz_regfile_17__15_), .A2(n6706), .ZN(n867) );
  NAND2_X2 U1571 ( .A1(regBoiz_regfile_17__14_), .A2(n6705), .ZN(n868) );
  NAND2_X2 U1573 ( .A1(regBoiz_regfile_17__13_), .A2(n6706), .ZN(n869) );
  NAND2_X2 U1575 ( .A1(regBoiz_regfile_17__12_), .A2(n6706), .ZN(n870) );
  NAND2_X2 U1577 ( .A1(regBoiz_regfile_17__11_), .A2(n841), .ZN(n871) );
  NAND2_X2 U1579 ( .A1(regBoiz_regfile_17__10_), .A2(n6706), .ZN(n872) );
  NAND2_X2 U1581 ( .A1(regBoiz_regfile_17__0_), .A2(n841), .ZN(n873) );
  NAND2_X2 U1582 ( .A1(n807), .A2(n99), .ZN(n841) );
  NAND2_X2 U1584 ( .A1(regBoiz_regfile_16__9_), .A2(n6702), .ZN(n875) );
  NAND2_X2 U1586 ( .A1(regBoiz_regfile_16__8_), .A2(n6701), .ZN(n876) );
  NAND2_X2 U1588 ( .A1(regBoiz_regfile_16__7_), .A2(n6700), .ZN(n877) );
  NAND2_X2 U1590 ( .A1(regBoiz_regfile_16__6_), .A2(n6701), .ZN(n878) );
  NAND2_X2 U1592 ( .A1(regBoiz_regfile_16__5_), .A2(n6700), .ZN(n879) );
  NAND2_X2 U1594 ( .A1(regBoiz_regfile_16__4_), .A2(n6701), .ZN(n880) );
  NAND2_X2 U1596 ( .A1(regBoiz_regfile_16__3_), .A2(n6700), .ZN(n881) );
  NAND2_X2 U1598 ( .A1(regBoiz_regfile_16__31_), .A2(n6701), .ZN(n882) );
  NAND2_X2 U1600 ( .A1(regBoiz_regfile_16__30_), .A2(n6702), .ZN(n883) );
  NAND2_X2 U1602 ( .A1(regBoiz_regfile_16__2_), .A2(n6702), .ZN(n884) );
  NAND2_X2 U1604 ( .A1(regBoiz_regfile_16__29_), .A2(n6702), .ZN(n885) );
  NAND2_X2 U1606 ( .A1(regBoiz_regfile_16__28_), .A2(n6702), .ZN(n886) );
  NAND2_X2 U1608 ( .A1(regBoiz_regfile_16__27_), .A2(n6702), .ZN(n887) );
  NAND2_X2 U1610 ( .A1(regBoiz_regfile_16__26_), .A2(n6702), .ZN(n888) );
  NAND2_X2 U1612 ( .A1(regBoiz_regfile_16__25_), .A2(n6702), .ZN(n889) );
  NAND2_X2 U1614 ( .A1(regBoiz_regfile_16__24_), .A2(n6702), .ZN(n890) );
  NAND2_X2 U1616 ( .A1(regBoiz_regfile_16__23_), .A2(n6702), .ZN(n891) );
  NAND2_X2 U1618 ( .A1(regBoiz_regfile_16__22_), .A2(n6702), .ZN(n892) );
  NAND2_X2 U1620 ( .A1(regBoiz_regfile_16__21_), .A2(n6702), .ZN(n893) );
  NAND2_X2 U1622 ( .A1(regBoiz_regfile_16__20_), .A2(n6702), .ZN(n894) );
  NAND2_X2 U1624 ( .A1(regBoiz_regfile_16__1_), .A2(n6702), .ZN(n895) );
  NAND2_X2 U1626 ( .A1(regBoiz_regfile_16__19_), .A2(n6702), .ZN(n896) );
  NAND2_X2 U1628 ( .A1(regBoiz_regfile_16__18_), .A2(n6702), .ZN(n897) );
  NAND2_X2 U1630 ( .A1(regBoiz_regfile_16__17_), .A2(n6702), .ZN(n898) );
  NAND2_X2 U1632 ( .A1(regBoiz_regfile_16__16_), .A2(n6702), .ZN(n899) );
  NAND2_X2 U1634 ( .A1(regBoiz_regfile_16__15_), .A2(n6702), .ZN(n900) );
  NAND2_X2 U1636 ( .A1(regBoiz_regfile_16__14_), .A2(n6702), .ZN(n901) );
  NAND2_X2 U1638 ( .A1(regBoiz_regfile_16__13_), .A2(n6702), .ZN(n902) );
  NAND2_X2 U1640 ( .A1(regBoiz_regfile_16__12_), .A2(n6702), .ZN(n903) );
  NAND2_X2 U1642 ( .A1(regBoiz_regfile_16__11_), .A2(n6702), .ZN(n904) );
  NAND2_X2 U1644 ( .A1(regBoiz_regfile_16__10_), .A2(n6702), .ZN(n905) );
  NAND2_X2 U1646 ( .A1(regBoiz_regfile_16__0_), .A2(n6702), .ZN(n906) );
  AND2_X2 U1648 ( .A1(n607), .A2(n907), .ZN(n807) );
  AND2_X2 U1649 ( .A1(wbRwh[4]), .A2(wbRegWrh), .ZN(n607) );
  NAND2_X2 U1651 ( .A1(regBoiz_regfile_15__9_), .A2(n6699), .ZN(n909) );
  NAND2_X2 U1659 ( .A1(regBoiz_regfile_15__5_), .A2(n6698), .ZN(n913) );
  NAND2_X2 U1661 ( .A1(regBoiz_regfile_15__4_), .A2(n6698), .ZN(n914) );
  NAND2_X2 U1663 ( .A1(regBoiz_regfile_15__3_), .A2(n6697), .ZN(n915) );
  NAND2_X2 U1665 ( .A1(regBoiz_regfile_15__31_), .A2(n6699), .ZN(n916) );
  NAND2_X2 U1667 ( .A1(regBoiz_regfile_15__30_), .A2(n6699), .ZN(n917) );
  NAND2_X2 U1669 ( .A1(regBoiz_regfile_15__2_), .A2(n6697), .ZN(n918) );
  NAND2_X2 U1671 ( .A1(regBoiz_regfile_15__29_), .A2(n6699), .ZN(n919) );
  NAND2_X2 U1673 ( .A1(regBoiz_regfile_15__28_), .A2(n6699), .ZN(n920) );
  NAND2_X2 U1675 ( .A1(regBoiz_regfile_15__27_), .A2(n6698), .ZN(n921) );
  NAND2_X2 U1677 ( .A1(regBoiz_regfile_15__26_), .A2(n6697), .ZN(n922) );
  NAND2_X2 U1679 ( .A1(regBoiz_regfile_15__25_), .A2(n908), .ZN(n923) );
  NAND2_X2 U1681 ( .A1(regBoiz_regfile_15__24_), .A2(n908), .ZN(n924) );
  NAND2_X2 U1685 ( .A1(regBoiz_regfile_15__22_), .A2(n908), .ZN(n926) );
  NAND2_X2 U1687 ( .A1(regBoiz_regfile_15__21_), .A2(n908), .ZN(n927) );
  NAND2_X2 U1689 ( .A1(regBoiz_regfile_15__20_), .A2(n908), .ZN(n928) );
  NAND2_X2 U1691 ( .A1(regBoiz_regfile_15__1_), .A2(n908), .ZN(n929) );
  NAND2_X2 U1693 ( .A1(regBoiz_regfile_15__19_), .A2(n908), .ZN(n930) );
  NAND2_X2 U1695 ( .A1(regBoiz_regfile_15__18_), .A2(n6699), .ZN(n931) );
  NAND2_X2 U1697 ( .A1(regBoiz_regfile_15__17_), .A2(n908), .ZN(n932) );
  NAND2_X2 U1701 ( .A1(regBoiz_regfile_15__15_), .A2(n6699), .ZN(n934) );
  NAND2_X2 U1703 ( .A1(regBoiz_regfile_15__14_), .A2(n908), .ZN(n935) );
  NAND2_X2 U1705 ( .A1(regBoiz_regfile_15__13_), .A2(n6699), .ZN(n936) );
  NAND2_X2 U1707 ( .A1(regBoiz_regfile_15__12_), .A2(n6699), .ZN(n937) );
  NAND2_X2 U1709 ( .A1(regBoiz_regfile_15__11_), .A2(n908), .ZN(n938) );
  NAND2_X2 U1713 ( .A1(regBoiz_regfile_15__0_), .A2(n908), .ZN(n940) );
  NAND2_X2 U1714 ( .A1(n941), .A2(n168), .ZN(n908) );
  NAND2_X2 U1716 ( .A1(regBoiz_regfile_14__9_), .A2(n6693), .ZN(n943) );
  NAND2_X2 U1718 ( .A1(regBoiz_regfile_14__8_), .A2(n6694), .ZN(n944) );
  NAND2_X2 U1722 ( .A1(regBoiz_regfile_14__6_), .A2(n6694), .ZN(n946) );
  NAND2_X2 U1724 ( .A1(regBoiz_regfile_14__5_), .A2(n6694), .ZN(n947) );
  NAND2_X2 U1728 ( .A1(regBoiz_regfile_14__3_), .A2(n6694), .ZN(n949) );
  NAND2_X2 U1730 ( .A1(regBoiz_regfile_14__31_), .A2(n6694), .ZN(n950) );
  NAND2_X2 U1732 ( .A1(regBoiz_regfile_14__30_), .A2(n6695), .ZN(n951) );
  NAND2_X2 U1734 ( .A1(regBoiz_regfile_14__2_), .A2(n6695), .ZN(n952) );
  NAND2_X2 U1736 ( .A1(regBoiz_regfile_14__29_), .A2(n6695), .ZN(n953) );
  NAND2_X2 U1738 ( .A1(regBoiz_regfile_14__28_), .A2(n6695), .ZN(n954) );
  NAND2_X2 U1742 ( .A1(regBoiz_regfile_14__26_), .A2(n6695), .ZN(n956) );
  NAND2_X2 U1744 ( .A1(regBoiz_regfile_14__25_), .A2(n6695), .ZN(n957) );
  NAND2_X2 U1746 ( .A1(regBoiz_regfile_14__24_), .A2(n6695), .ZN(n958) );
  NAND2_X2 U1748 ( .A1(regBoiz_regfile_14__23_), .A2(n6695), .ZN(n959) );
  NAND2_X2 U1750 ( .A1(regBoiz_regfile_14__22_), .A2(n6695), .ZN(n960) );
  NAND2_X2 U1752 ( .A1(regBoiz_regfile_14__21_), .A2(n6695), .ZN(n961) );
  NAND2_X2 U1754 ( .A1(regBoiz_regfile_14__20_), .A2(n6695), .ZN(n962) );
  NAND2_X2 U1756 ( .A1(regBoiz_regfile_14__1_), .A2(n6695), .ZN(n963) );
  NAND2_X2 U1758 ( .A1(regBoiz_regfile_14__19_), .A2(n6695), .ZN(n964) );
  NAND2_X2 U1760 ( .A1(regBoiz_regfile_14__18_), .A2(n6695), .ZN(n965) );
  NAND2_X2 U1762 ( .A1(regBoiz_regfile_14__17_), .A2(n6695), .ZN(n966) );
  NAND2_X2 U1766 ( .A1(regBoiz_regfile_14__15_), .A2(n6694), .ZN(n968) );
  NAND2_X2 U1768 ( .A1(regBoiz_regfile_14__14_), .A2(n6695), .ZN(n969) );
  NAND2_X2 U1770 ( .A1(regBoiz_regfile_14__13_), .A2(n6695), .ZN(n970) );
  NAND2_X2 U1772 ( .A1(regBoiz_regfile_14__12_), .A2(n6695), .ZN(n971) );
  NAND2_X2 U1774 ( .A1(regBoiz_regfile_14__11_), .A2(n6695), .ZN(n972) );
  NAND2_X2 U1776 ( .A1(regBoiz_regfile_14__10_), .A2(n6695), .ZN(n973) );
  NAND2_X2 U1778 ( .A1(regBoiz_regfile_14__0_), .A2(n6695), .ZN(n974) );
  NAND2_X2 U1779 ( .A1(n941), .A2(n203), .ZN(n942) );
  NAND2_X2 U1781 ( .A1(regBoiz_regfile_13__9_), .A2(n6691), .ZN(n976) );
  NAND2_X2 U1783 ( .A1(regBoiz_regfile_13__8_), .A2(n6689), .ZN(n977) );
  NAND2_X2 U1787 ( .A1(regBoiz_regfile_13__6_), .A2(n6690), .ZN(n979) );
  NAND2_X2 U1789 ( .A1(regBoiz_regfile_13__5_), .A2(n6689), .ZN(n980) );
  NAND2_X2 U1793 ( .A1(regBoiz_regfile_13__3_), .A2(n6690), .ZN(n982) );
  NAND2_X2 U1795 ( .A1(regBoiz_regfile_13__31_), .A2(n6689), .ZN(n983) );
  NAND2_X2 U1797 ( .A1(regBoiz_regfile_13__30_), .A2(n6691), .ZN(n984) );
  NAND2_X2 U1799 ( .A1(regBoiz_regfile_13__2_), .A2(n6691), .ZN(n985) );
  NAND2_X2 U1801 ( .A1(regBoiz_regfile_13__29_), .A2(n6691), .ZN(n986) );
  NAND2_X2 U1803 ( .A1(regBoiz_regfile_13__28_), .A2(n6691), .ZN(n987) );
  NAND2_X2 U1805 ( .A1(regBoiz_regfile_13__27_), .A2(n6691), .ZN(n988) );
  NAND2_X2 U1807 ( .A1(regBoiz_regfile_13__26_), .A2(n6691), .ZN(n989) );
  NAND2_X2 U1809 ( .A1(regBoiz_regfile_13__25_), .A2(n6691), .ZN(n990) );
  NAND2_X2 U1811 ( .A1(regBoiz_regfile_13__24_), .A2(n6691), .ZN(n991) );
  NAND2_X2 U1813 ( .A1(regBoiz_regfile_13__23_), .A2(n6691), .ZN(n992) );
  NAND2_X2 U1815 ( .A1(regBoiz_regfile_13__22_), .A2(n6691), .ZN(n993) );
  NAND2_X2 U1817 ( .A1(regBoiz_regfile_13__21_), .A2(n6691), .ZN(n994) );
  NAND2_X2 U1819 ( .A1(regBoiz_regfile_13__20_), .A2(n6691), .ZN(n995) );
  NAND2_X2 U1821 ( .A1(regBoiz_regfile_13__1_), .A2(n6691), .ZN(n996) );
  NAND2_X2 U1823 ( .A1(regBoiz_regfile_13__19_), .A2(n6691), .ZN(n997) );
  NAND2_X2 U1825 ( .A1(regBoiz_regfile_13__18_), .A2(n6691), .ZN(n998) );
  NAND2_X2 U1827 ( .A1(regBoiz_regfile_13__17_), .A2(n6691), .ZN(n999) );
  NAND2_X2 U1829 ( .A1(regBoiz_regfile_13__16_), .A2(n6691), .ZN(n1000) );
  NAND2_X2 U1831 ( .A1(regBoiz_regfile_13__15_), .A2(n6691), .ZN(n1001) );
  NAND2_X2 U1833 ( .A1(regBoiz_regfile_13__14_), .A2(n6691), .ZN(n1002) );
  NAND2_X2 U1835 ( .A1(regBoiz_regfile_13__13_), .A2(n6691), .ZN(n1003) );
  NAND2_X2 U1837 ( .A1(regBoiz_regfile_13__12_), .A2(n6691), .ZN(n1004) );
  NAND2_X2 U1839 ( .A1(regBoiz_regfile_13__11_), .A2(n6691), .ZN(n1005) );
  NAND2_X2 U1841 ( .A1(regBoiz_regfile_13__10_), .A2(n6691), .ZN(n1006) );
  NAND2_X2 U1843 ( .A1(regBoiz_regfile_13__0_), .A2(n6691), .ZN(n1007) );
  NAND2_X2 U1847 ( .A1(regBoiz_regfile_12__9_), .A2(n6688), .ZN(n1010) );
  NAND2_X2 U1849 ( .A1(regBoiz_regfile_12__8_), .A2(n6687), .ZN(n1011) );
  NAND2_X2 U1851 ( .A1(regBoiz_regfile_12__7_), .A2(n6686), .ZN(n1012) );
  NAND2_X2 U1853 ( .A1(regBoiz_regfile_12__6_), .A2(n6687), .ZN(n1013) );
  NAND2_X2 U1855 ( .A1(regBoiz_regfile_12__5_), .A2(n6686), .ZN(n1014) );
  NAND2_X2 U1857 ( .A1(regBoiz_regfile_12__4_), .A2(n6686), .ZN(n1015) );
  NAND2_X2 U1859 ( .A1(regBoiz_regfile_12__3_), .A2(n6687), .ZN(n1016) );
  NAND2_X2 U1861 ( .A1(regBoiz_regfile_12__31_), .A2(n6686), .ZN(n1017) );
  NAND2_X2 U1863 ( .A1(regBoiz_regfile_12__30_), .A2(n6688), .ZN(n1018) );
  NAND2_X2 U1865 ( .A1(regBoiz_regfile_12__2_), .A2(n6688), .ZN(n1019) );
  NAND2_X2 U1867 ( .A1(regBoiz_regfile_12__29_), .A2(n6688), .ZN(n1020) );
  NAND2_X2 U1869 ( .A1(regBoiz_regfile_12__28_), .A2(n6688), .ZN(n1021) );
  NAND2_X2 U1871 ( .A1(regBoiz_regfile_12__27_), .A2(n6688), .ZN(n1022) );
  NAND2_X2 U1873 ( .A1(regBoiz_regfile_12__26_), .A2(n6688), .ZN(n1023) );
  NAND2_X2 U1875 ( .A1(regBoiz_regfile_12__25_), .A2(n6688), .ZN(n1024) );
  NAND2_X2 U1877 ( .A1(regBoiz_regfile_12__24_), .A2(n6688), .ZN(n1025) );
  NAND2_X2 U1879 ( .A1(regBoiz_regfile_12__23_), .A2(n6688), .ZN(n1026) );
  NAND2_X2 U1881 ( .A1(regBoiz_regfile_12__22_), .A2(n6688), .ZN(n1027) );
  NAND2_X2 U1883 ( .A1(regBoiz_regfile_12__21_), .A2(n6688), .ZN(n1028) );
  NAND2_X2 U1885 ( .A1(regBoiz_regfile_12__20_), .A2(n6688), .ZN(n1029) );
  NAND2_X2 U1887 ( .A1(regBoiz_regfile_12__1_), .A2(n6688), .ZN(n1030) );
  NAND2_X2 U1889 ( .A1(regBoiz_regfile_12__19_), .A2(n6688), .ZN(n1031) );
  NAND2_X2 U1891 ( .A1(regBoiz_regfile_12__18_), .A2(n6688), .ZN(n1032) );
  NAND2_X2 U1893 ( .A1(regBoiz_regfile_12__17_), .A2(n6688), .ZN(n1033) );
  NAND2_X2 U1895 ( .A1(regBoiz_regfile_12__16_), .A2(n6688), .ZN(n1034) );
  NAND2_X2 U1897 ( .A1(regBoiz_regfile_12__15_), .A2(n6688), .ZN(n1035) );
  NAND2_X2 U1899 ( .A1(regBoiz_regfile_12__14_), .A2(n6688), .ZN(n1036) );
  NAND2_X2 U1901 ( .A1(regBoiz_regfile_12__13_), .A2(n6688), .ZN(n1037) );
  NAND2_X2 U1903 ( .A1(regBoiz_regfile_12__12_), .A2(n6688), .ZN(n1038) );
  NAND2_X2 U1905 ( .A1(regBoiz_regfile_12__11_), .A2(n6688), .ZN(n1039) );
  NAND2_X2 U1907 ( .A1(regBoiz_regfile_12__10_), .A2(n6688), .ZN(n1040) );
  NAND2_X2 U1909 ( .A1(regBoiz_regfile_12__0_), .A2(n6688), .ZN(n1041) );
  AND2_X2 U1911 ( .A1(wbRwh[2]), .A2(n1042), .ZN(n941) );
  NAND2_X2 U1913 ( .A1(regBoiz_regfile_11__9_), .A2(n6685), .ZN(n1044) );
  NAND2_X2 U1915 ( .A1(regBoiz_regfile_11__8_), .A2(n6683), .ZN(n1045) );
  NAND2_X2 U1917 ( .A1(regBoiz_regfile_11__7_), .A2(n6683), .ZN(n1046) );
  NAND2_X2 U1919 ( .A1(regBoiz_regfile_11__6_), .A2(n6684), .ZN(n1047) );
  NAND2_X2 U1921 ( .A1(regBoiz_regfile_11__5_), .A2(n6683), .ZN(n1048) );
  NAND2_X2 U1923 ( .A1(regBoiz_regfile_11__4_), .A2(n6684), .ZN(n1049) );
  NAND2_X2 U1925 ( .A1(regBoiz_regfile_11__3_), .A2(n6684), .ZN(n1050) );
  NAND2_X2 U1927 ( .A1(regBoiz_regfile_11__31_), .A2(n6685), .ZN(n1051) );
  NAND2_X2 U1929 ( .A1(regBoiz_regfile_11__30_), .A2(n6685), .ZN(n1052) );
  NAND2_X2 U1931 ( .A1(regBoiz_regfile_11__2_), .A2(n6685), .ZN(n1053) );
  NAND2_X2 U1933 ( .A1(regBoiz_regfile_11__29_), .A2(n6685), .ZN(n1054) );
  NAND2_X2 U1935 ( .A1(regBoiz_regfile_11__28_), .A2(n6685), .ZN(n1055) );
  NAND2_X2 U1937 ( .A1(regBoiz_regfile_11__27_), .A2(n6685), .ZN(n1056) );
  NAND2_X2 U1939 ( .A1(regBoiz_regfile_11__26_), .A2(n6685), .ZN(n1057) );
  NAND2_X2 U1941 ( .A1(regBoiz_regfile_11__25_), .A2(n6685), .ZN(n1058) );
  NAND2_X2 U1943 ( .A1(regBoiz_regfile_11__24_), .A2(n6685), .ZN(n1059) );
  NAND2_X2 U1945 ( .A1(regBoiz_regfile_11__23_), .A2(n6685), .ZN(n1060) );
  NAND2_X2 U1947 ( .A1(regBoiz_regfile_11__22_), .A2(n6685), .ZN(n1061) );
  NAND2_X2 U1949 ( .A1(regBoiz_regfile_11__21_), .A2(n6685), .ZN(n1062) );
  NAND2_X2 U1951 ( .A1(regBoiz_regfile_11__20_), .A2(n6685), .ZN(n1063) );
  NAND2_X2 U1953 ( .A1(regBoiz_regfile_11__1_), .A2(n6685), .ZN(n1064) );
  NAND2_X2 U1955 ( .A1(regBoiz_regfile_11__19_), .A2(n6685), .ZN(n1065) );
  NAND2_X2 U1957 ( .A1(regBoiz_regfile_11__18_), .A2(n6685), .ZN(n1066) );
  NAND2_X2 U1959 ( .A1(regBoiz_regfile_11__17_), .A2(n6685), .ZN(n1067) );
  NAND2_X2 U1961 ( .A1(regBoiz_regfile_11__16_), .A2(n6683), .ZN(n1068) );
  NAND2_X2 U1963 ( .A1(regBoiz_regfile_11__15_), .A2(n6685), .ZN(n1069) );
  NAND2_X2 U1965 ( .A1(regBoiz_regfile_11__14_), .A2(n6685), .ZN(n1070) );
  NAND2_X2 U1967 ( .A1(regBoiz_regfile_11__13_), .A2(n6684), .ZN(n1071) );
  NAND2_X2 U1969 ( .A1(regBoiz_regfile_11__12_), .A2(n6685), .ZN(n1072) );
  NAND2_X2 U1971 ( .A1(regBoiz_regfile_11__11_), .A2(n6685), .ZN(n1073) );
  NAND2_X2 U1973 ( .A1(regBoiz_regfile_11__10_), .A2(n6685), .ZN(n1074) );
  NAND2_X2 U1975 ( .A1(regBoiz_regfile_11__0_), .A2(n6685), .ZN(n1075) );
  NAND2_X2 U1976 ( .A1(n168), .A2(n100), .ZN(n1043) );
  AND2_X2 U1977 ( .A1(wbRwh[1]), .A2(wbRwh[0]), .ZN(n168) );
  NAND2_X2 U1979 ( .A1(regBoiz_regfile_10__9_), .A2(net367597), .ZN(n1077) );
  NAND2_X2 U1981 ( .A1(regBoiz_regfile_10__8_), .A2(net367595), .ZN(n1078) );
  NAND2_X2 U1983 ( .A1(regBoiz_regfile_10__7_), .A2(net367593), .ZN(n1079) );
  NAND2_X2 U1985 ( .A1(regBoiz_regfile_10__6_), .A2(net367595), .ZN(n1080) );
  NAND2_X2 U1987 ( .A1(regBoiz_regfile_10__5_), .A2(net367593), .ZN(n1081) );
  NAND2_X2 U1989 ( .A1(regBoiz_regfile_10__4_), .A2(net367593), .ZN(n1082) );
  NAND2_X2 U1991 ( .A1(regBoiz_regfile_10__3_), .A2(net367595), .ZN(n1083) );
  NAND2_X2 U1995 ( .A1(regBoiz_regfile_10__30_), .A2(net367597), .ZN(n1085) );
  NAND2_X2 U1997 ( .A1(regBoiz_regfile_10__2_), .A2(net367597), .ZN(n1086) );
  NAND2_X2 U1999 ( .A1(regBoiz_regfile_10__29_), .A2(net367597), .ZN(n1087) );
  NAND2_X2 U2001 ( .A1(regBoiz_regfile_10__28_), .A2(net367597), .ZN(n1088) );
  NAND2_X2 U2005 ( .A1(regBoiz_regfile_10__26_), .A2(net367597), .ZN(n1090) );
  NAND2_X2 U2007 ( .A1(regBoiz_regfile_10__25_), .A2(net367597), .ZN(n1091) );
  NAND2_X2 U2009 ( .A1(regBoiz_regfile_10__24_), .A2(net367597), .ZN(n1092) );
  NAND2_X2 U2011 ( .A1(regBoiz_regfile_10__23_), .A2(net367597), .ZN(n1093) );
  NAND2_X2 U2013 ( .A1(regBoiz_regfile_10__22_), .A2(net367597), .ZN(n1094) );
  NAND2_X2 U2015 ( .A1(regBoiz_regfile_10__21_), .A2(net367597), .ZN(n1095) );
  NAND2_X2 U2017 ( .A1(regBoiz_regfile_10__20_), .A2(net367597), .ZN(n1096) );
  NAND2_X2 U2019 ( .A1(regBoiz_regfile_10__1_), .A2(net367597), .ZN(n1097) );
  NAND2_X2 U2021 ( .A1(regBoiz_regfile_10__19_), .A2(net367597), .ZN(n1098) );
  NAND2_X2 U2023 ( .A1(regBoiz_regfile_10__18_), .A2(net367597), .ZN(n1099) );
  NAND2_X2 U2025 ( .A1(regBoiz_regfile_10__17_), .A2(net367597), .ZN(n1100) );
  NAND2_X2 U2027 ( .A1(regBoiz_regfile_10__16_), .A2(net367597), .ZN(n1101) );
  NAND2_X2 U2029 ( .A1(regBoiz_regfile_10__15_), .A2(net367597), .ZN(n1102) );
  NAND2_X2 U2031 ( .A1(regBoiz_regfile_10__14_), .A2(net367597), .ZN(n1103) );
  NAND2_X2 U2033 ( .A1(regBoiz_regfile_10__13_), .A2(net367597), .ZN(n1104) );
  NAND2_X2 U2035 ( .A1(regBoiz_regfile_10__12_), .A2(net367597), .ZN(n1105) );
  NAND2_X2 U2037 ( .A1(regBoiz_regfile_10__11_), .A2(net367597), .ZN(n1106) );
  NAND2_X2 U2039 ( .A1(regBoiz_regfile_10__10_), .A2(net367597), .ZN(n1107) );
  NAND2_X2 U2041 ( .A1(regBoiz_regfile_10__0_), .A2(net367597), .ZN(n1108) );
  AND2_X2 U2043 ( .A1(n1042), .A2(n5482), .ZN(n100) );
  AND2_X2 U2045 ( .A1(wbRwh[3]), .A2(n271), .ZN(n1042) );
  AND2_X2 U2046 ( .A1(wbRwh[1]), .A2(n5511), .ZN(n203) );
  NAND2_X2 U2049 ( .A1(regBoiz_regfile_0__9_), .A2(n6680), .ZN(n1110) );
  NAND2_X2 U2052 ( .A1(regBoiz_regfile_0__8_), .A2(n6678), .ZN(n1111) );
  NAND2_X2 U2055 ( .A1(regBoiz_regfile_0__7_), .A2(n6679), .ZN(n1112) );
  NAND2_X2 U2058 ( .A1(regBoiz_regfile_0__6_), .A2(n6678), .ZN(n1113) );
  NAND2_X2 U2061 ( .A1(regBoiz_regfile_0__5_), .A2(n6679), .ZN(n1114) );
  NAND2_X2 U2064 ( .A1(regBoiz_regfile_0__4_), .A2(n6678), .ZN(n1115) );
  NAND2_X2 U2067 ( .A1(regBoiz_regfile_0__3_), .A2(n6679), .ZN(n1116) );
  NAND2_X2 U2070 ( .A1(regBoiz_regfile_0__31_), .A2(n6680), .ZN(n1117) );
  NAND2_X2 U2073 ( .A1(regBoiz_regfile_0__30_), .A2(n6680), .ZN(n1118) );
  NAND2_X2 U2076 ( .A1(regBoiz_regfile_0__2_), .A2(n6680), .ZN(n1119) );
  NAND2_X2 U2079 ( .A1(regBoiz_regfile_0__29_), .A2(n6680), .ZN(n1120) );
  NAND2_X2 U2082 ( .A1(regBoiz_regfile_0__28_), .A2(n6680), .ZN(n1121) );
  NAND2_X2 U2085 ( .A1(regBoiz_regfile_0__27_), .A2(n6680), .ZN(n1122) );
  NAND2_X2 U2088 ( .A1(regBoiz_regfile_0__26_), .A2(n6680), .ZN(n1123) );
  NAND2_X2 U2091 ( .A1(regBoiz_regfile_0__25_), .A2(n6680), .ZN(n1124) );
  NAND2_X2 U2094 ( .A1(regBoiz_regfile_0__24_), .A2(n6680), .ZN(n1125) );
  NAND2_X2 U2097 ( .A1(regBoiz_regfile_0__23_), .A2(n6680), .ZN(n1126) );
  NAND2_X2 U2100 ( .A1(regBoiz_regfile_0__22_), .A2(n6680), .ZN(n1127) );
  NAND2_X2 U2103 ( .A1(regBoiz_regfile_0__21_), .A2(n6680), .ZN(n1128) );
  NAND2_X2 U2106 ( .A1(regBoiz_regfile_0__20_), .A2(n6680), .ZN(n1129) );
  NAND2_X2 U2109 ( .A1(regBoiz_regfile_0__1_), .A2(n6680), .ZN(n1130) );
  NAND2_X2 U2112 ( .A1(regBoiz_regfile_0__19_), .A2(n6680), .ZN(n1131) );
  NAND2_X2 U2115 ( .A1(regBoiz_regfile_0__18_), .A2(n6680), .ZN(n1132) );
  NAND2_X2 U2118 ( .A1(regBoiz_regfile_0__17_), .A2(n6680), .ZN(n1133) );
  NAND2_X2 U2121 ( .A1(regBoiz_regfile_0__16_), .A2(n6680), .ZN(n1134) );
  NAND2_X2 U2124 ( .A1(regBoiz_regfile_0__15_), .A2(n6679), .ZN(n1135) );
  NAND2_X2 U2127 ( .A1(regBoiz_regfile_0__14_), .A2(n6680), .ZN(n1136) );
  NAND2_X2 U2130 ( .A1(regBoiz_regfile_0__13_), .A2(n6678), .ZN(n1137) );
  NAND2_X2 U2133 ( .A1(regBoiz_regfile_0__12_), .A2(n6680), .ZN(n1138) );
  NAND2_X2 U2136 ( .A1(regBoiz_regfile_0__11_), .A2(n6680), .ZN(n1139) );
  NAND2_X2 U2139 ( .A1(regBoiz_regfile_0__10_), .A2(n6680), .ZN(n1140) );
  NAND2_X2 U2142 ( .A1(regBoiz_regfile_0__0_), .A2(n6680), .ZN(n1141) );
  NAND2_X2 U2143 ( .A1(n305), .A2(n134), .ZN(n1109) );
  AND2_X2 U2145 ( .A1(n907), .A2(n271), .ZN(n305) );
  AOI22_X2 U2151 ( .A1(n1146), .A2(daddr[3]), .B1(drData[3]), .B2(n1147), .ZN(
        n1145) );
  AOI22_X2 U2153 ( .A1(n1146), .A2(daddr[2]), .B1(drData[2]), .B2(n1147), .ZN(
        n1149) );
  AOI22_X2 U2155 ( .A1(n1146), .A2(daddr[1]), .B1(drData[1]), .B2(n1147), .ZN(
        n1151) );
  AOI22_X2 U2157 ( .A1(n1146), .A2(daddr[0]), .B1(drData[0]), .B2(n1147), .ZN(
        n1153) );
  OAI221_X2 U2158 ( .B1(n5328), .B2(n13712), .C1(n5689), .C2(n5377), .A(n1157), 
        .ZN(n3498) );
  OAI221_X2 U2160 ( .B1(n5321), .B2(n13712), .C1(n5689), .C2(n5376), .A(n1162), 
        .ZN(n3531) );
  OAI221_X2 U2163 ( .B1(n5327), .B2(n13712), .C1(n5689), .C2(n5375), .A(n1165), 
        .ZN(n3564) );
  OAI221_X2 U2166 ( .B1(n5320), .B2(n13712), .C1(n5689), .C2(n5374), .A(n1168), 
        .ZN(n3597) );
  OAI221_X2 U2169 ( .B1(n5379), .B2(n13712), .C1(n5689), .C2(n5330), .A(n1171), 
        .ZN(n3630) );
  OAI221_X2 U2172 ( .B1(n5378), .B2(n13712), .C1(n5689), .C2(n5329), .A(n1174), 
        .ZN(n3663) );
  OAI221_X2 U2175 ( .B1(n5326), .B2(n13712), .C1(n5689), .C2(n5373), .A(n1177), 
        .ZN(n3696) );
  OAI221_X2 U2178 ( .B1(n5325), .B2(n13712), .C1(n5689), .C2(n5372), .A(n1180), 
        .ZN(n3729) );
  OAI221_X2 U2181 ( .B1(n5324), .B2(n13712), .C1(n5689), .C2(n5371), .A(n1183), 
        .ZN(n3762) );
  OAI221_X2 U2184 ( .B1(n5503), .B2(n13712), .C1(n5689), .C2(n5370), .A(n1186), 
        .ZN(n3795) );
  OAI221_X2 U2187 ( .B1(n5502), .B2(n13712), .C1(n5689), .C2(n5369), .A(n1189), 
        .ZN(n3828) );
  OAI221_X2 U2190 ( .B1(n5501), .B2(n13712), .C1(n5689), .C2(n5368), .A(n1192), 
        .ZN(n3861) );
  OAI221_X2 U2193 ( .B1(n5323), .B2(n13712), .C1(n5689), .C2(n5367), .A(n1195), 
        .ZN(n3894) );
  OAI221_X2 U2196 ( .B1(n5500), .B2(n13712), .C1(n5689), .C2(n5366), .A(n1198), 
        .ZN(n3927) );
  OAI221_X2 U2199 ( .B1(n5499), .B2(n13712), .C1(n5689), .C2(n5365), .A(n1201), 
        .ZN(n3960) );
  OAI221_X2 U2202 ( .B1(n5322), .B2(n13712), .C1(n5689), .C2(n5364), .A(n1204), 
        .ZN(n3993) );
  OAI211_X2 U2205 ( .C1(n1206), .C2(n1207), .A(n1147), .B(n6943), .ZN(n1205)
         );
  AND3_X2 U2206 ( .A1(drData[15]), .A2(aluDExtOp), .A3(n1208), .ZN(n1207) );
  OAI221_X2 U2209 ( .B1(n1210), .B2(n6959), .C1(n13676), .C2(n1213), .A(n1214), 
        .ZN(n4026) );
  AOI22_X2 U2211 ( .A1(n1146), .A2(daddr[15]), .B1(aluPC8[15]), .B2(aluJAL), 
        .ZN(n1210) );
  OAI211_X2 U2212 ( .C1(n5498), .C2(n13712), .A(n1214), .B(n1216), .ZN(n4059)
         );
  AOI22_X2 U2213 ( .A1(drData[14]), .A2(n13674), .B1(aluPC8[14]), .B2(aluJAL), 
        .ZN(n1216) );
  OAI211_X2 U2215 ( .C1(n5488), .C2(n13712), .A(n1214), .B(n1219), .ZN(n4092)
         );
  AOI22_X2 U2216 ( .A1(drData[13]), .A2(n13674), .B1(aluPC8[13]), .B2(aluJAL), 
        .ZN(n1219) );
  OAI211_X2 U2218 ( .C1(n5491), .C2(n13712), .A(n1214), .B(n1221), .ZN(n4125)
         );
  AOI22_X2 U2219 ( .A1(drData[12]), .A2(n13674), .B1(aluPC8[12]), .B2(aluJAL), 
        .ZN(n1221) );
  OAI211_X2 U2221 ( .C1(n5497), .C2(n13712), .A(n1214), .B(n1223), .ZN(n4158)
         );
  AOI22_X2 U2222 ( .A1(drData[11]), .A2(n13674), .B1(aluPC8[11]), .B2(aluJAL), 
        .ZN(n1223) );
  OAI211_X2 U2224 ( .C1(n5496), .C2(n13712), .A(n1214), .B(n1225), .ZN(n4191)
         );
  AOI22_X2 U2225 ( .A1(drData[10]), .A2(n13674), .B1(aluPC8[10]), .B2(aluJAL), 
        .ZN(n1225) );
  OAI211_X2 U2227 ( .C1(n5495), .C2(n13712), .A(n1214), .B(n1227), .ZN(n4224)
         );
  AOI22_X2 U2228 ( .A1(drData[9]), .A2(n13674), .B1(aluPC8[9]), .B2(aluJAL), 
        .ZN(n1227) );
  OAI211_X2 U2230 ( .C1(n5487), .C2(n13712), .A(n1214), .B(n1229), .ZN(n4257)
         );
  AOI22_X2 U2231 ( .A1(drData[8]), .A2(n13674), .B1(aluPC8[8]), .B2(aluJAL), 
        .ZN(n1229) );
  OAI211_X2 U2233 ( .C1(n1209), .C2(n1208), .A(n1147), .B(n6943), .ZN(n1213)
         );
  NAND2_X2 U2236 ( .A1(n1206), .A2(n1147), .ZN(n1214) );
  AND3_X2 U2237 ( .A1(aluDExtOp), .A2(n5318), .A3(drData[7]), .ZN(n1206) );
  AOI22_X2 U2243 ( .A1(n1146), .A2(daddr[6]), .B1(drData[6]), .B2(n1147), .ZN(
        n1234) );
  AOI22_X2 U2245 ( .A1(n1146), .A2(daddr[5]), .B1(drData[5]), .B2(n1147), .ZN(
        n1236) );
  AOI22_X2 U2247 ( .A1(n1146), .A2(daddr[4]), .B1(drData[4]), .B2(n1147), .ZN(
        n1238) );
  NAND2_X2 U2485 ( .A1(pcIn[9]), .A2(n6960), .ZN(n3446) );
  OR2_X2 U2486 ( .A1(pcRst), .A2(pcIn[9]), .ZN(n3447) );
  NAND2_X2 U2495 ( .A1(pcIn[8]), .A2(n6960), .ZN(n3448) );
  OR2_X2 U2496 ( .A1(pcRst), .A2(pcIn[8]), .ZN(n3449) );
  NAND2_X2 U2506 ( .A1(pcIn[7]), .A2(n6960), .ZN(n3450) );
  OR2_X2 U2507 ( .A1(pcRst), .A2(pcIn[7]), .ZN(n3451) );
  NAND2_X2 U2516 ( .A1(pcIn[6]), .A2(n6960), .ZN(n3452) );
  OR2_X2 U2517 ( .A1(pcRst), .A2(pcIn[6]), .ZN(n3453) );
  NAND2_X2 U2524 ( .A1(pcIn[5]), .A2(n6960), .ZN(n3454) );
  OR2_X2 U2525 ( .A1(pcRst), .A2(pcIn[5]), .ZN(n3455) );
  NAND2_X2 U2533 ( .A1(pcIn[4]), .A2(n6960), .ZN(n3456) );
  OR2_X2 U2534 ( .A1(pcRst), .A2(pcIn[4]), .ZN(n3457) );
  NAND2_X2 U2541 ( .A1(pcIn[3]), .A2(n6960), .ZN(n3458) );
  OR2_X2 U2542 ( .A1(pcRst), .A2(pcIn[3]), .ZN(n3459) );
  NAND2_X2 U2557 ( .A1(pcIn[31]), .A2(n6960), .ZN(n3402) );
  OR2_X2 U2558 ( .A1(pcRst), .A2(pcIn[31]), .ZN(n3403) );
  NAND2_X2 U2584 ( .A1(pcIn[30]), .A2(n6960), .ZN(n3404) );
  OR2_X2 U2585 ( .A1(pcRst), .A2(pcIn[30]), .ZN(n3405) );
  NAND2_X2 U2590 ( .A1(pcIn[2]), .A2(n6960), .ZN(n3460) );
  OR2_X2 U2591 ( .A1(pcRst), .A2(pcIn[2]), .ZN(n3461) );
  NAND2_X2 U2606 ( .A1(pcIn[29]), .A2(n6960), .ZN(n3406) );
  OR2_X2 U2607 ( .A1(pcRst), .A2(pcIn[29]), .ZN(n3407) );
  NAND2_X2 U2625 ( .A1(pcIn[28]), .A2(n6961), .ZN(n3408) );
  OR2_X2 U2626 ( .A1(pcRst), .A2(pcIn[28]), .ZN(n3409) );
  NAND2_X2 U2640 ( .A1(pcIn[27]), .A2(n6961), .ZN(n3410) );
  OR2_X2 U2641 ( .A1(pcRst), .A2(pcIn[27]), .ZN(n3411) );
  NAND2_X2 U2655 ( .A1(pcIn[26]), .A2(n6961), .ZN(n3412) );
  OR2_X2 U2656 ( .A1(pcRst), .A2(pcIn[26]), .ZN(n3413) );
  NAND2_X2 U2672 ( .A1(pcIn[25]), .A2(n6961), .ZN(n3414) );
  OR2_X2 U2673 ( .A1(pcRst), .A2(pcIn[25]), .ZN(n3415) );
  NAND2_X2 U2688 ( .A1(pcIn[24]), .A2(n6961), .ZN(n3416) );
  OR2_X2 U2689 ( .A1(pcRst), .A2(pcIn[24]), .ZN(n3417) );
  NAND2_X2 U2704 ( .A1(pcIn[23]), .A2(n6961), .ZN(n3418) );
  OR2_X2 U2705 ( .A1(pcRst), .A2(pcIn[23]), .ZN(n3419) );
  NAND2_X2 U2720 ( .A1(pcIn[22]), .A2(n6961), .ZN(n3420) );
  OR2_X2 U2721 ( .A1(pcRst), .A2(pcIn[22]), .ZN(n3421) );
  NAND2_X2 U2736 ( .A1(pcIn[21]), .A2(n6961), .ZN(n3422) );
  OR2_X2 U2737 ( .A1(pcRst), .A2(pcIn[21]), .ZN(n3423) );
  NAND2_X2 U2752 ( .A1(pcIn[20]), .A2(n6961), .ZN(n3424) );
  OR2_X2 U2753 ( .A1(pcRst), .A2(pcIn[20]), .ZN(n3425) );
  NAND2_X2 U2759 ( .A1(pcIn[1]), .A2(n6961), .ZN(n3462) );
  OR2_X2 U2760 ( .A1(pcRst), .A2(pcIn[1]), .ZN(n3463) );
  NAND2_X2 U2775 ( .A1(pcIn[19]), .A2(n6961), .ZN(n3426) );
  OR2_X2 U2776 ( .A1(pcRst), .A2(pcIn[19]), .ZN(n3427) );
  NAND2_X2 U2791 ( .A1(pcIn[18]), .A2(n6960), .ZN(n3428) );
  OR2_X2 U2792 ( .A1(pcRst), .A2(pcIn[18]), .ZN(n3429) );
  NAND2_X2 U2807 ( .A1(pcIn[17]), .A2(n6961), .ZN(n3430) );
  OR2_X2 U2808 ( .A1(pcRst), .A2(pcIn[17]), .ZN(n3431) );
  NAND2_X2 U2823 ( .A1(pcIn[16]), .A2(n6960), .ZN(n3432) );
  OR2_X2 U2824 ( .A1(pcRst), .A2(pcIn[16]), .ZN(n3433) );
  NAND2_X2 U2838 ( .A1(pcIn[15]), .A2(n6961), .ZN(n3434) );
  OR2_X2 U2839 ( .A1(pcRst), .A2(pcIn[15]), .ZN(n3435) );
  NAND2_X2 U2853 ( .A1(pcIn[14]), .A2(n6960), .ZN(n3436) );
  OR2_X2 U2854 ( .A1(pcRst), .A2(pcIn[14]), .ZN(n3437) );
  NAND2_X2 U2868 ( .A1(pcIn[13]), .A2(n6961), .ZN(n3438) );
  OR2_X2 U2869 ( .A1(pcRst), .A2(pcIn[13]), .ZN(n3439) );
  NAND2_X2 U2883 ( .A1(pcIn[12]), .A2(n6960), .ZN(n3440) );
  OR2_X2 U2884 ( .A1(pcRst), .A2(pcIn[12]), .ZN(n3441) );
  NAND2_X2 U2897 ( .A1(pcIn[11]), .A2(n6961), .ZN(n3442) );
  OR2_X2 U2898 ( .A1(pcRst), .A2(pcIn[11]), .ZN(n3443) );
  NAND2_X2 U2962 ( .A1(pcIn[10]), .A2(n6960), .ZN(n3444) );
  OR2_X2 U2963 ( .A1(pcRst), .A2(pcIn[10]), .ZN(n3445) );
  NAND2_X2 U2978 ( .A1(pcIn[0]), .A2(n6961), .ZN(n3464) );
  OR2_X2 U2980 ( .A1(pcRst), .A2(pcIn[0]), .ZN(n3465) );
  OR4_X2 U3136 ( .A1(ifInst[21]), .A2(ifInst[22]), .A3(ifInst[20]), .A4(n2010), 
        .ZN(n2009) );
  NOR4_X2 U3144 ( .A1(n2014), .A2(ifInst[14]), .A3(ifInst[16]), .A4(ifInst[15]), .ZN(n2013) );
  OR3_X2 U3145 ( .A1(ifInst[18]), .A2(ifInst[19]), .A3(ifInst[17]), .ZN(n2014)
         );
  XNOR2_X2 U3227 ( .A(ifInst[27]), .B(ifInst[28]), .ZN(n2082) );
  OR4_X2 U3329 ( .A1(net368481), .A2(aluBoi_multBoi_count_0_), .A3(
        aluBoi_multBoi_count_1_), .A4(aluBoi_multBoi_count_2_), .ZN(n2105) );
  NAND2_X2 U3515 ( .A1(n2202), .A2(net100619), .ZN(aluBoi_multBoi_N73) );
  XNOR2_X2 U3516 ( .A(aluBoi_multBoi_count_2_), .B(n2203), .ZN(n2202) );
  NAND2_X2 U3518 ( .A1(n2204), .A2(net100619), .ZN(aluBoi_multBoi_N72) );
  XOR2_X2 U3519 ( .A(aluBoi_multBoi_count_1_), .B(aluBoi_multBoi_count_0_), 
        .Z(n2204) );
  NAND2_X2 U3520 ( .A1(aluBoi_multBoi_count_0_), .A2(net100619), .ZN(
        aluBoi_multBoi_N71) );
  OAI22_X2 U4197 ( .A1(idOut_18_), .A2(n5716), .B1(n13538), .B2(n5391), .ZN(
        n2842) );
  AOI22_X2 U4199 ( .A1(n2844), .A2(n2847), .B1(n13538), .B2(n5391), .ZN(n2840)
         );
  NAND2_X2 U4252 ( .A1(idOut_19_), .A2(idOut_20_), .ZN(aluBoi_condBoi_N24) );
  OAI22_X2 U4255 ( .A1(n5371), .A2(n6611), .B1(n6607), .B2(n5636), .ZN(n4530)
         );
  OAI22_X2 U4258 ( .A1(n5370), .A2(n6611), .B1(n6607), .B2(n5635), .ZN(n4531)
         );
  OAI22_X2 U4261 ( .A1(n5369), .A2(n6611), .B1(n6607), .B2(n5634), .ZN(n4532)
         );
  OAI22_X2 U4264 ( .A1(n5368), .A2(n6611), .B1(n6607), .B2(n5633), .ZN(n4533)
         );
  OAI22_X2 U4267 ( .A1(n5367), .A2(n6611), .B1(n6607), .B2(n5632), .ZN(n4534)
         );
  OAI22_X2 U4270 ( .A1(n5366), .A2(n6611), .B1(n6607), .B2(n5631), .ZN(n4535)
         );
  OAI22_X2 U4273 ( .A1(n5365), .A2(n6611), .B1(n6607), .B2(n5630), .ZN(n4536)
         );
  OAI22_X2 U4276 ( .A1(n5364), .A2(n6611), .B1(n6607), .B2(n5629), .ZN(n4537)
         );
  AOI22_X2 U4280 ( .A1(aluPC8[15]), .A2(n6609), .B1(n6608), .B2(idOut_54_), 
        .ZN(n2983) );
  AOI22_X2 U4282 ( .A1(aluPC8[14]), .A2(n6609), .B1(n6608), .B2(idOut_53_), 
        .ZN(n2984) );
  AOI22_X2 U4286 ( .A1(aluPC8[13]), .A2(n6609), .B1(n6608), .B2(idOut_52_), 
        .ZN(n2986) );
  AOI22_X2 U4288 ( .A1(aluPC8[12]), .A2(n6609), .B1(n6608), .B2(idOut_51_), 
        .ZN(n2987) );
  AOI22_X2 U4290 ( .A1(aluPC8[11]), .A2(n6609), .B1(n6608), .B2(idOut_50_), 
        .ZN(n2988) );
  AOI22_X2 U4292 ( .A1(aluPC8[10]), .A2(n6609), .B1(n6608), .B2(idOut_49_), 
        .ZN(n2989) );
  AOI22_X2 U4294 ( .A1(aluPC8[9]), .A2(n6609), .B1(n6608), .B2(idOut_48_), 
        .ZN(n2990) );
  AOI22_X2 U4296 ( .A1(aluPC8[8]), .A2(n6609), .B1(n6608), .B2(idOut_47_), 
        .ZN(n2991) );
  AOI22_X2 U4298 ( .A1(aluPC8[7]), .A2(n6609), .B1(n6608), .B2(idOut_46_), 
        .ZN(n2992) );
  OAI22_X2 U4299 ( .A1(n5358), .A2(n6611), .B1(n6607), .B2(n5628), .ZN(n4547)
         );
  OAI22_X2 U4302 ( .A1(n5357), .A2(n6611), .B1(n6607), .B2(n5627), .ZN(n4548)
         );
  OAI22_X2 U4305 ( .A1(n5356), .A2(n6611), .B1(n6607), .B2(n5626), .ZN(n4549)
         );
  OAI22_X2 U4310 ( .A1(n5362), .A2(n6611), .B1(n6607), .B2(n5625), .ZN(n4550)
         );
  OAI22_X2 U4313 ( .A1(n5361), .A2(n6611), .B1(n6607), .B2(n5624), .ZN(n4551)
         );
  OAI22_X2 U4316 ( .A1(n5360), .A2(n6611), .B1(n6607), .B2(n5623), .ZN(n4552)
         );
  OAI22_X2 U4319 ( .A1(n5359), .A2(n6611), .B1(n6607), .B2(n5622), .ZN(n4553)
         );
  AOI22_X2 U4427 ( .A1(n6609), .A2(dWr), .B1(n6608), .B2(idOut_34_), .ZN(n3083) );
  OAI22_X2 U4594 ( .A1(n5384), .A2(n6611), .B1(n6607), .B2(n5621), .ZN(n4718)
         );
  OAI22_X2 U4738 ( .A1(n5353), .A2(n6611), .B1(n6607), .B2(n5620), .ZN(n4794)
         );
  OAI211_X2 U4842 ( .C1(n5595), .C2(n3353), .A(n3354), .B(n3355), .ZN(n4801)
         );
  OAI211_X2 U4845 ( .C1(n5594), .C2(n3353), .A(n3354), .B(n3357), .ZN(n4796)
         );
  AOI22_X2 U4846 ( .A1(n3356), .A2(n6832), .B1(aluRw[3]), .B2(n6609), .ZN(
        n3357) );
  OAI211_X2 U4848 ( .C1(n5593), .C2(n3353), .A(n3354), .B(n3358), .ZN(n4800)
         );
  AOI22_X2 U4849 ( .A1(n3356), .A2(n6823), .B1(aluRw[2]), .B2(n6609), .ZN(
        n3358) );
  OAI211_X2 U4851 ( .C1(n5592), .C2(n3353), .A(n3354), .B(n3359), .ZN(n4797)
         );
  AOI22_X2 U4852 ( .A1(n3356), .A2(n6804), .B1(aluRw[1]), .B2(n6609), .ZN(
        n3359) );
  OAI22_X2 U4854 ( .A1(n5318), .A2(n6611), .B1(n6607), .B2(n5619), .ZN(n4716)
         );
  OAI211_X2 U4857 ( .C1(n5591), .C2(n3353), .A(n3354), .B(n3360), .ZN(n4798)
         );
  AOI22_X2 U4858 ( .A1(n3356), .A2(net369154), .B1(n5898), .B2(n6609), .ZN(
        n3360) );
  NAND2_X2 U4860 ( .A1(idOut_38_), .A2(n6608), .ZN(n3353) );
  NAND2_X2 U4881 ( .A1(idOut_26_), .A2(n6608), .ZN(n3354) );
  OAI22_X2 U4903 ( .A1(n5519), .A2(n6611), .B1(n6607), .B2(n5583), .ZN(n4714)
         );
  OAI22_X2 U4928 ( .A1(n5377), .A2(n6611), .B1(n6607), .B2(n5618), .ZN(n4522)
         );
  OAI22_X2 U4931 ( .A1(n5376), .A2(n6611), .B1(n6607), .B2(n5617), .ZN(n4523)
         );
  OAI22_X2 U4934 ( .A1(n5375), .A2(n6611), .B1(n6607), .B2(n5616), .ZN(n4524)
         );
  OAI22_X2 U4937 ( .A1(n5374), .A2(n6611), .B1(n6607), .B2(n5615), .ZN(n4525)
         );
  OAI22_X2 U4940 ( .A1(n5330), .A2(n6611), .B1(n6607), .B2(n5614), .ZN(n4526)
         );
  OAI22_X2 U4943 ( .A1(n5329), .A2(n6611), .B1(n6607), .B2(n5613), .ZN(n4527)
         );
  OAI22_X2 U4946 ( .A1(n5373), .A2(n6611), .B1(n6607), .B2(n5612), .ZN(n4528)
         );
  OAI22_X2 U4949 ( .A1(n5372), .A2(n6611), .B1(n6607), .B2(n5611), .ZN(n4529)
         );
  AOI22_X2 U4955 ( .A1(n6609), .A2(aluRegWrOut), .B1(n6608), .B2(idRegWr), 
        .ZN(n3391) );
  DFFR_X2 ifBoi_reglol_60__regBoi_curData_reg ( .D(n13604), .CK(clk), .RN(
        n6916), .Q(ifInst[28]) );
  DFFR_X2 ifBoi_reglol_59__regBoi_curData_reg ( .D(n13603), .CK(clk), .RN(
        n6915), .Q(ifInst[27]) );
  DFFR_X2 ifBoi_reglol_32__regBoi_curData_reg ( .D(n13576), .CK(clk), .RN(
        n6897), .Q(idBoi_temPC_0_), .QN(n5459) );
  DFFR_X2 idBoi_reggal_76__regBoi_curData_reg ( .D(n13613), .CK(clk), .RN(
        n6894), .Q(regBoiz_N15), .QN(net369138) );
  DFFR_X2 aluBoi_aluReg_2__regBoi_curData_reg ( .D(n4799), .CK(clk), .RN(n6886), .Q(aluJAL), .QN(n5689) );
  DFFR_X2 idBoi_reggal_37__regBoi_curData_reg ( .D(n4787), .CK(clk), .RN(n6881), .QN(n5714) );
  DFFR_X2 idBoi_reggal_81__regBoi_curData_reg ( .D(n13618), .CK(clk), .RN(
        n6895), .Q(net368800), .QN(net368712) );
  DFFR_X2 idBoi_reggal_83__regBoi_curData_reg ( .D(n13620), .CK(clk), .RN(
        n6895), .Q(regBoiz_N12), .QN(net375279) );
  DFFR_X2 idBoi_reggal_84__regBoi_curData_reg ( .D(n13621), .CK(clk), .RN(
        n6878), .Q(net375642), .QN(net368681) );
  DFFR_X2 idBoi_reggal_85__regBoi_curData_reg ( .D(n13622), .CK(clk), .RN(
        n6895), .Q(n6370), .QN(n6413) );
  DFFR_X2 idBoi_reggal_82__regBoi_curData_reg ( .D(n13619), .CK(clk), .RN(
        n6879), .Q(net375527), .QN(net368676) );
  DFFR_X2 regBoiz_regfile_reg_21__4_ ( .D(n3619), .CK(clk), .RN(n6855), .Q(
        regBoiz_regfile_21__4_), .QN(n6505) );
  DFFR_X2 regBoiz_regfile_reg_29__4_ ( .D(n3627), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_29__4_), .QN(n6504) );
  DFFR_X2 regBoiz_regfile_reg_23__9_ ( .D(n3786), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__9_), .QN(n6502) );
  DFFR_X2 regBoiz_regfile_reg_31__9_ ( .D(n3794), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__9_), .QN(n6501) );
  DFFR_X2 regBoiz_regfile_reg_23__3_ ( .D(n3588), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__3_), .QN(n6497) );
  DFFR_X2 regBoiz_regfile_reg_31__3_ ( .D(n3596), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__3_), .QN(n6496) );
  DFFR_X2 regBoiz_regfile_reg_19__4_ ( .D(n3617), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__4_), .QN(n6491) );
  DFFR_X2 regBoiz_regfile_reg_27__4_ ( .D(n3625), .CK(clk), .RN(n6847), .Q(
        regBoiz_regfile_27__4_), .QN(n6490) );
  DFFR_X2 regBoiz_regfile_reg_23__4_ ( .D(n3621), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__4_), .QN(n6488) );
  DFFR_X2 regBoiz_regfile_reg_31__4_ ( .D(n3629), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__4_), .QN(n6487) );
  DFFR_X2 regBoiz_regfile_reg_19__9_ ( .D(n3782), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_19__9_), .QN(n6485) );
  DFFR_X2 regBoiz_regfile_reg_27__9_ ( .D(n3790), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_27__9_), .QN(n6484) );
  DFFR_X2 regBoiz_regfile_reg_22__4_ ( .D(n3620), .CK(clk), .RN(n6853), .Q(
        regBoiz_regfile_22__4_), .QN(n6482) );
  DFFR_X2 regBoiz_regfile_reg_30__4_ ( .D(n3628), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_30__4_), .QN(n6481) );
  DFFR_X2 regBoiz_regfile_reg_22__9_ ( .D(n3785), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_22__9_), .QN(n6479) );
  DFFR_X2 regBoiz_regfile_reg_30__9_ ( .D(n3793), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__9_), .QN(n6478) );
  DFFR_X2 regBoiz_regfile_reg_30__10_ ( .D(n3826), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__10_), .QN(n6472) );
  DFFR_X2 regBoiz_regfile_reg_31__10_ ( .D(n3827), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_31__10_), .QN(n6471) );
  DFFR_X2 regBoiz_regfile_reg_15__4_ ( .D(n3613), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__4_), .QN(n6469) );
  DFFR_X2 regBoiz_regfile_reg_29__9_ ( .D(n3792), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__9_), .QN(n6467) );
  DFFR_X2 regBoiz_regfile_reg_15__9_ ( .D(n3778), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__9_), .QN(n6465) );
  DFFR_X2 regBoiz_regfile_reg_30__3_ ( .D(n3595), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__3_), .QN(n6463) );
  DFFR_X2 regBoiz_regfile_reg_29__3_ ( .D(n3594), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__3_), .QN(n6462) );
  DFFR_X2 regBoiz_regfile_reg_27__3_ ( .D(n3592), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_27__3_), .QN(n6460) );
  DFFR_X2 regBoiz_regfile_reg_14__3_ ( .D(n3579), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__3_), .QN(n6459) );
  DFFR_X2 regBoiz_regfile_reg_15__3_ ( .D(n3580), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__3_), .QN(n6458) );
  DFFR_X2 regBoiz_regfile_reg_15__10_ ( .D(n3811), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_15__10_), .QN(n6446) );
  DFFR_X2 regBoiz_regfile_reg_28__4_ ( .D(n3626), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_28__4_), .QN(n6443) );
  DFFR_X2 regBoiz_regfile_reg_28__9_ ( .D(n3791), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_28__9_), .QN(n6348) );
  DFFR_X2 regBoiz_regfile_reg_29__10_ ( .D(n3825), .CK(clk), .RN(n6929), .Q(
        regBoiz_regfile_29__10_), .QN(n6455) );
  DFFR_X2 regBoiz_regfile_reg_15__7_ ( .D(n3712), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__7_), .QN(n6454) );
  DFFR_X2 regBoiz_regfile_reg_27__10_ ( .D(n3823), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__10_), .QN(n6452) );
  DFFR_X2 regBoiz_regfile_reg_23__10_ ( .D(n3819), .CK(clk), .RN(n6921), .Q(
        regBoiz_regfile_23__10_), .QN(n6450) );
  DFFR_X2 regBoiz_regfile_reg_26__9_ ( .D(n3789), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__9_), .QN(n6448) );
  DFFR_X2 regBoiz_regfile_reg_11__4_ ( .D(n3609), .CK(clk), .RN(n6869), .Q(
        regBoiz_regfile_11__4_), .QN(net368926) );
  DFFR_X2 regBoiz_regfile_reg_7__4_ ( .D(n3605), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_7__4_), .QN(n6340) );
  DFFR_X2 regBoiz_regfile_reg_26__4_ ( .D(n3624), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__4_), .QN(n6353) );
  DFFR_X2 regBoiz_regfile_reg_14__9_ ( .D(n3777), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__9_), .QN(n6444) );
  DFFR_X2 regBoiz_regfile_reg_14__4_ ( .D(n3612), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_14__4_), .QN(n6338) );
  DFFR_X2 regBoiz_regfile_reg_25__4_ ( .D(n3623), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_25__4_), .QN(n6341) );
  DFFR_X2 regBoiz_regfile_reg_21__9_ ( .D(n3784), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_21__9_) );
  DFFR_X2 regBoiz_regfile_reg_13__9_ ( .D(n3776), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_13__9_) );
  DFFR_X2 regBoiz_regfile_reg_9__9_ ( .D(n3772), .CK(clk), .RN(n6943), .Q(
        regBoiz_regfile_9__9_), .QN(n6406) );
  DFFR_X2 regBoiz_regfile_reg_7__9_ ( .D(n3770), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__9_) );
  DFFR_X2 regBoiz_regfile_reg_3__10_ ( .D(n3799), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__10_), .QN(n6405) );
  DFFR_X2 regBoiz_regfile_reg_11__10_ ( .D(n3807), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_11__10_), .QN(n6404) );
  DFFR_X2 regBoiz_regfile_reg_26__10_ ( .D(n3822), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_26__10_) );
  DFFR_X2 regBoiz_regfile_reg_22__10_ ( .D(n3818), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__10_) );
  DFFR_X2 regBoiz_regfile_reg_28__10_ ( .D(n3824), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__10_) );
  DFFR_X2 regBoiz_regfile_reg_21__10_ ( .D(n3817), .CK(clk), .RN(n6919), .Q(
        regBoiz_regfile_21__10_), .QN(n6329) );
  DFFR_X2 regBoiz_regfile_reg_14__10_ ( .D(n3810), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__10_), .QN(n6395) );
  DFFR_X2 aluBoi_aluReg_44__regBoi_curData_reg ( .D(n4781), .CK(clk), .RN(
        n6885), .Q(daddr[0]), .QN(net375393) );
  DFFR_X2 regBoiz_regfile_reg_19__10_ ( .D(n3815), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__10_) );
  DFFR_X2 regBoiz_regfile_reg_25__10_ ( .D(n3821), .CK(clk), .RN(n6924), .Q(
        regBoiz_regfile_25__10_) );
  DFFR_X2 regBoiz_regfile_reg_10__28_ ( .D(n4400), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__28_), .QN(n6391) );
  DFFR_X2 regBoiz_regfile_reg_26__28_ ( .D(n4416), .CK(clk), .RN(n6848), .Q(
        regBoiz_regfile_26__28_), .QN(n6390) );
  DFFR_X2 regBoiz_regfile_reg_22__23_ ( .D(n4247), .CK(clk), .RN(n6920), .Q(
        regBoiz_regfile_22__23_), .QN(n6383) );
  DFFR_X2 regBoiz_regfile_reg_30__23_ ( .D(n4255), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__23_), .QN(n6382) );
  DFFR_X2 regBoiz_regfile_reg_31__23_ ( .D(n4256), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__23_), .QN(n6377) );
  DFFR_X2 regBoiz_regfile_reg_23__23_ ( .D(n4248), .CK(clk), .RN(n6922), .Q(
        regBoiz_regfile_23__23_) );
  DFFR_X2 regBoiz_regfile_reg_30__13_ ( .D(n3925), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__13_), .QN(net375528) );
  DFFR_X2 regBoiz_regfile_reg_28__13_ ( .D(n3923), .CK(clk), .RN(n6846), .Q(
        regBoiz_regfile_28__13_), .QN(net375526) );
  DFFR_X2 regBoiz_regfile_reg_10__31_ ( .D(n4499), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__31_), .QN(n6292) );
  DFFR_X2 regBoiz_regfile_reg_16__27_ ( .D(n4373), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__27_) );
  DFFR_X2 regBoiz_regfile_reg_24__27_ ( .D(n4381), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__27_) );
  DFFR_X2 regBoiz_regfile_reg_18__23_ ( .D(n4243), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__23_), .QN(n6364) );
  DFFR_X2 regBoiz_regfile_reg_26__23_ ( .D(n4251), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__23_), .QN(n6363) );
  DFFR_X2 regBoiz_regfile_reg_20__9_ ( .D(n3783), .CK(clk), .RN(n6918), .Q(
        regBoiz_regfile_20__9_), .QN(n6347) );
  DFFR_X2 regBoiz_regfile_reg_13__4_ ( .D(n3611), .CK(clk), .RN(n6867), .Q(
        regBoiz_regfile_13__4_), .QN(n6336) );
  DFFR_X2 regBoiz_regfile_reg_31__2_ ( .D(n3563), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__2_), .QN(n6310) );
  DFFR_X2 regBoiz_regfile_reg_31__1_ ( .D(n3530), .CK(clk), .RN(n6934), .Q(
        regBoiz_regfile_31__1_), .QN(n6332) );
  DFFR_X2 regBoiz_regfile_reg_20__4_ ( .D(n3618), .CK(clk), .RN(n6856), .Q(
        regBoiz_regfile_20__4_), .QN(n6326) );
  DFFR_X2 regBoiz_regfile_reg_6__4_ ( .D(n3604), .CK(clk), .RN(n6836), .Q(
        regBoiz_regfile_6__4_), .QN(n6304) );
  DFFR_X2 regBoiz_regfile_reg_14__7_ ( .D(n3711), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__7_), .QN(n6281) );
  DFFR_X2 regBoiz_regfile_reg_11__7_ ( .D(n3708), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__7_), .QN(n6323) );
  DFFR_X2 regBoiz_regfile_reg_13__7_ ( .D(n3710), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_13__7_), .QN(n6308) );
  DFFR_X2 regBoiz_regfile_reg_31__8_ ( .D(n3761), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__8_), .QN(n6321) );
  DFFR_X2 regBoiz_regfile_reg_12__4_ ( .D(n3610), .CK(clk), .RN(n6868), .Q(
        regBoiz_regfile_12__4_), .QN(n6319) );
  DFFR_X2 regBoiz_regfile_reg_10__4_ ( .D(n3608), .CK(clk), .RN(n6871), .Q(
        regBoiz_regfile_10__4_), .QN(n6317) );
  DFFR_X2 regBoiz_regfile_reg_17__4_ ( .D(n3615), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_17__4_), .QN(n6303) );
  DFFR_X2 regBoiz_regfile_reg_15__8_ ( .D(n3745), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__8_) );
  DFFR_X2 regBoiz_regfile_reg_9__4_ ( .D(n3607), .CK(clk), .RN(n6937), .Q(
        regBoiz_regfile_9__4_), .QN(n6314) );
  DFFR_X2 regBoiz_regfile_reg_3__4_ ( .D(n3601), .CK(clk), .RN(n6840), .Q(
        regBoiz_regfile_3__4_), .QN(net375768) );
  DFFR_X2 regBoiz_regfile_reg_5__4_ ( .D(n3603), .CK(clk), .RN(n6837), .Q(
        regBoiz_regfile_5__4_), .QN(n6312) );
  DFFR_X2 regBoiz_regfile_reg_30__1_ ( .D(n3529), .CK(clk), .RN(n6932), .Q(
        regBoiz_regfile_30__1_), .QN(n6298) );
  DFFR_X2 regBoiz_regfile_reg_7__7_ ( .D(n3704), .CK(clk), .RN(n6941), .Q(
        regBoiz_regfile_7__7_), .QN(n6306) );
  DFFR_X2 regBoiz_regfile_reg_7__1_ ( .D(n3506), .CK(clk), .RN(n6940), .Q(
        regBoiz_regfile_7__1_) );
  DFFR_X2 regBoiz_regfile_reg_28__1_ ( .D(n3527), .CK(clk), .RN(n6928), .Q(
        regBoiz_regfile_28__1_), .QN(n6297) );
  DFFR_X2 regBoiz_regfile_reg_29__1_ ( .D(n3528), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__1_), .QN(n6296) );
  DFF_X1 aluBoi_multBoi_runProd_reg_60_ ( .D(aluBoi_multBoi_N66), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[56]), .QN(n5572) );
  DFFR_X2 regBoiz_regfile_reg_25__9_ ( .D(n3788), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_25__9_), .QN(n6233) );
  DFFR_X2 regBoiz_regfile_reg_2__31_ ( .D(n4491), .CK(clk), .RN(n6844), .Q(
        regBoiz_regfile_2__31_), .QN(n6291) );
  DFFR_X2 regBoiz_regfile_reg_30__29_ ( .D(n4453), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_30__29_), .QN(n6283) );
  DFFR_X2 regBoiz_regfile_reg_31__13_ ( .D(n3926), .CK(clk), .RN(n6842), .Q(
        regBoiz_regfile_31__13_) );
  DFFR_X2 regBoiz_regfile_reg_19__28_ ( .D(n4409), .CK(clk), .RN(n6859), .Q(
        regBoiz_regfile_19__28_) );
  DFFR_X2 regBoiz_regfile_reg_31__6_ ( .D(n3695), .CK(clk), .RN(n6841), .Q(
        regBoiz_regfile_31__6_) );
  DFFR_X2 regBoiz_regfile_reg_15__6_ ( .D(n3679), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__6_) );
  DFFR_X2 regBoiz_regfile_reg_18__28_ ( .D(n4408), .CK(clk), .RN(n6860), .Q(
        regBoiz_regfile_18__28_) );
  DFFR_X2 regBoiz_regfile_reg_15__23_ ( .D(n4240), .CK(clk), .RN(n6910), .Q(
        regBoiz_regfile_15__23_) );
  DFFR_X2 regBoiz_regfile_reg_27__23_ ( .D(n4252), .CK(clk), .RN(n6927), .Q(
        regBoiz_regfile_27__23_) );
  DFFR_X2 aluBoi_aluReg_40__regBoi_curData_reg ( .D(n4797), .CK(clk), .RN(
        n6885), .Q(aluRw[1]), .QN(n4995) );
  DFFR_X2 regBoiz_regfile_reg_14__16_ ( .D(n4008), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__16_), .QN(n5247) );
  DFFR_X2 regBoiz_regfile_reg_14__29_ ( .D(n4437), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__29_), .QN(n6171) );
  DFFR_X2 aluBoi_aluReg_39__regBoi_curData_reg ( .D(n4798), .CK(clk), .RN(
        n6885), .Q(aluRw[0]), .QN(n5897) );
  DFFR_X2 regBoiz_regfile_reg_26__29_ ( .D(n4449), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__29_), .QN(n6175) );
  DFFR_X2 regBoiz_regfile_reg_24__23_ ( .D(n4249), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__23_) );
  DFFR_X2 aluBoi_aluReg_42__regBoi_curData_reg ( .D(n4796), .CK(clk), .RN(
        n6885), .Q(aluRw[3]), .QN(n5949) );
  DFF_X1 aluBoi_multBoi_runProd_reg_45_ ( .D(aluBoi_multBoi_N51), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[41]), .QN(net376800) );
  DFFR_X2 regBoiz_regfile_reg_15__16_ ( .D(n4009), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_15__16_) );
  DFFR_X2 regBoiz_regfile_reg_8__31_ ( .D(n4497), .CK(clk), .RN(n6904), .Q(
        regBoiz_regfile_8__31_) );
  DFFR_X2 regBoiz_regfile_reg_11__29_ ( .D(n4434), .CK(clk), .RN(n6905), .Q(
        regBoiz_regfile_11__29_), .QN(n6030) );
  DFFR_X2 regBoiz_regfile_reg_24__28_ ( .D(n4414), .CK(clk), .RN(n6851), .Q(
        regBoiz_regfile_24__28_) );
  DFF_X1 aluBoi_multBoi_runProd_reg_57_ ( .D(aluBoi_multBoi_N63), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[53]), .QN(n5521) );
  DFFR_X2 idBoi_reggal_2__regBoi_curData_reg ( .D(n4815), .CK(clk), .RN(n6881), 
        .Q(aluBoi_imm32w_2_), .QN(n6073) );
  DFFR_X2 regBoiz_regfile_reg_29__5_ ( .D(n3660), .CK(clk), .RN(n6930), .Q(
        regBoiz_regfile_29__5_), .QN(n6043) );
  DFF_X1 aluBoi_multBoi_runProd_reg_62_ ( .D(aluBoi_multBoi_N68), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[58]), .QN(n5558) );
  DFFR_X2 regBoiz_regfile_reg_3__12_ ( .D(n3865), .CK(clk), .RN(n6935), .Q(
        regBoiz_regfile_3__12_), .QN(n6025) );
  DFFR_X2 regBoiz_regfile_reg_1__12_ ( .D(n3863), .CK(clk), .RN(n6916), .Q(
        regBoiz_regfile_1__12_), .QN(n6024) );
  DFFR_X2 regBoiz_regfile_reg_31__16_ ( .D(n4025), .CK(clk), .RN(n6933), .Q(
        regBoiz_regfile_31__16_), .QN(n6021) );
  DFFR_X2 regBoiz_regfile_reg_15__12_ ( .D(n3877), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_15__12_) );
  DFFR_X2 regBoiz_regfile_reg_17__28_ ( .D(n4407), .CK(clk), .RN(n6862), .Q(
        regBoiz_regfile_17__28_), .QN(n6017) );
  DFFR_X2 ifBoi_reglol_34__regBoi_curData_reg ( .D(n13578), .CK(clk), .RN(
        n6897), .Q(idBoi_temPC_2_), .QN(n5312) );
  DFFR_X2 aluBoi_aluReg_43__regBoi_curData_reg ( .D(n4801), .CK(clk), .RN(
        n6889), .Q(aluRw[4]) );
  DFFR_X2 idBoi_reggal_1__regBoi_curData_reg ( .D(n4817), .CK(clk), .RN(n6939), 
        .Q(aluBoi_imm32w_1_), .QN(n5994) );
  DFFR_X2 regBoiz_regfile_reg_14__12_ ( .D(n3876), .CK(clk), .RN(n6908), .Q(
        regBoiz_regfile_14__12_) );
  DFFR_X2 regBoiz_regfile_reg_15__22_ ( .D(n4207), .CK(clk), .RN(n6865), .Q(
        regBoiz_regfile_15__22_) );
  DFFR_X2 regBoiz_regfile_reg_6__29_ ( .D(n4429), .CK(clk), .RN(n6939), .Q(
        regBoiz_regfile_6__29_) );
  DFFR_X1 ifBoi_reglol_33__regBoi_curData_reg ( .D(n13577), .CK(clk), .RN(
        n6877), .Q(idBoi_temPC_1_), .QN(n5940) );
  DFFR_X1 regBoiz_regfile_reg_15__26_ ( .D(n4339), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_15__26_), .QN(n5932) );
  NAND2_X2 U2003 ( .A1(regBoiz_regfile_10__27_), .A2(net367597), .ZN(n1089) );
  NAND2_X2 U628 ( .A1(regBoiz_regfile_2__27_), .A2(net367221), .ZN(n386) );
  DFFR_X2 regBoiz_regfile_reg_24__18_ ( .D(n4084), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__18_) );
  DFF_X1 aluBoi_multBoi_runProd_reg_56_ ( .D(aluBoi_multBoi_N62), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[52]), .QN(n5483) );
  DFFR_X2 regBoiz_regfile_reg_22__28_ ( .D(n4412), .CK(clk), .RN(n6854), .Q(
        regBoiz_regfile_22__28_) );
  DFFR_X2 idBoi_reggal_88__regBoi_curData_reg ( .D(n4701), .CK(clk), .RN(n6878), .Q(idOut_88_), .QN(n5725) );
  DFFR_X2 aluBoi_aluReg_71__regBoi_curData_reg ( .D(n4767), .CK(clk), .RN(
        n6884), .Q(daddr[27]), .QN(n5379) );
  DFFR_X2 idBoi_reggal_3__regBoi_curData_reg ( .D(n4831), .CK(clk), .RN(n6893), 
        .Q(aluBoi_imm32w_3_) );
  DFFR_X2 idBoi_reggal_0__regBoi_curData_reg ( .D(n4821), .CK(clk), .RN(n6883), 
        .Q(aluBoi_imm32w_0_) );
  DFFR_X2 aluBoi_aluReg_70__regBoi_curData_reg ( .D(n4769), .CK(clk), .RN(
        n6890), .Q(daddr[26]), .QN(n5378) );
  DFF_X1 aluBoi_multBoi_runProd_reg_44_ ( .D(aluBoi_multBoi_N50), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[40]), .QN(n5569) );
  DFFRS_X1 ifBoi_pcOut_reg_28_ ( .D(n4573), .CK(clk), .RN(n3409), .SN(n3408), 
        .Q(iaddr[28]) );
  DFF_X1 aluBoi_multBoi_runProd_reg_41_ ( .D(aluBoi_multBoi_N47), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[37]) );
  DFFR_X2 idBoi_reggal_4__regBoi_curData_reg ( .D(n4812), .CK(clk), .RN(n6880), 
        .Q(aluBoi_imm32w_4_) );
  DFF_X1 aluBoi_multBoi_runProd_reg_40_ ( .D(aluBoi_multBoi_N46), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[36]), .QN(n5687) );
  DFF_X1 aluBoi_multBoi_runProd_reg_47_ ( .D(n5049), .CK(clk), .Q(
        aluBoi_multBoi_temppp[43]), .QN(n5685) );
  DFF_X1 aluBoi_multBoi_runProd_reg_42_ ( .D(aluBoi_multBoi_N48), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[38]), .QN(n5681) );
  DFF_X1 aluBoi_multBoi_runProd_reg_37_ ( .D(aluBoi_multBoi_N43), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[33]), .QN(n5680) );
  DFFR_X2 idBoi_reggal_79__regBoi_curData_reg ( .D(n13616), .CK(clk), .RN(
        n6879), .Q(regBoiz_N18), .QN(n5677) );
  DFF_X1 aluBoi_multBoi_runProd_reg_50_ ( .D(aluBoi_multBoi_N56), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[46]), .QN(n5646) );
  DFF_X1 aluBoi_multBoi_runProd_reg_61_ ( .D(aluBoi_multBoi_N67), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[57]), .QN(n5348) );
  DFF_X1 aluBoi_multBoi_runProd_reg_39_ ( .D(aluBoi_multBoi_N45), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[35]), .QN(n5639) );
  DFF_X1 aluBoi_multBoi_runProd_reg_46_ ( .D(aluBoi_multBoi_N52), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[42]), .QN(n5596) );
  DFF_X1 aluBoi_multBoi_runProd_reg_43_ ( .D(aluBoi_multBoi_N49), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[39]), .QN(n5585) );
  DFFRS_X1 ifBoi_pcOut_reg_27_ ( .D(n4578), .CK(clk), .RN(n3411), .SN(n3410), 
        .Q(iaddr[27]), .QN(n5580) );
  DFF_X1 aluBoi_multBoi_runProd_reg_51_ ( .D(aluBoi_multBoi_N57), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[47]), .QN(n5573) );
  DFFRS_X1 ifBoi_pcOut_reg_29_ ( .D(n4568), .CK(clk), .RN(n3407), .SN(n3406), 
        .Q(iaddr[29]), .QN(n5571) );
  DFFRS_X1 ifBoi_pcOut_reg_21_ ( .D(n4608), .CK(clk), .RN(n3423), .SN(n3422), 
        .Q(iaddr[21]), .QN(n5562) );
  DFF_X1 aluBoi_multBoi_runProd_reg_49_ ( .D(aluBoi_multBoi_N55), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[45]), .QN(n5560) );
  DFFRS_X1 ifBoi_pcOut_reg_24_ ( .D(n4593), .CK(clk), .RN(n3417), .SN(n3416), 
        .Q(iaddr[24]), .QN(n5559) );
  DFF_X1 aluBoi_multBoi_runProd_reg_55_ ( .D(aluBoi_multBoi_N61), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[51]), .QN(n5551) );
  DFFR_X2 regBoiz_regfile_reg_17__21_ ( .D(n4176), .CK(clk), .RN(n6912), .Q(
        regBoiz_regfile_17__21_), .QN(n5545) );
  DFF_X1 aluBoi_multBoi_runProd_reg_59_ ( .D(aluBoi_multBoi_N65), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[55]), .QN(n5537) );
  DFFR_X2 regBoiz_regfile_reg_16__21_ ( .D(n4175), .CK(clk), .RN(n6911), .Q(
        regBoiz_regfile_16__21_), .QN(n5536) );
  DFFR_X2 regBoiz_regfile_reg_0__21_ ( .D(n4159), .CK(clk), .RN(n6902), .Q(
        regBoiz_regfile_0__21_), .QN(n5535) );
  DFFR_X2 regBoiz_regfile_reg_18__21_ ( .D(n4177), .CK(clk), .RN(n6914), .Q(
        regBoiz_regfile_18__21_), .QN(n5534) );
  DFFR_X2 regBoiz_regfile_reg_8__21_ ( .D(n4167), .CK(clk), .RN(n6942), .Q(
        regBoiz_regfile_8__21_), .QN(n5531) );
  DFFR_X2 regBoiz_regfile_reg_26__15_ ( .D(n3987), .CK(clk), .RN(n6849), .Q(
        regBoiz_regfile_26__15_), .QN(n5530) );
  DFFR_X2 regBoiz_regfile_reg_24__15_ ( .D(n3985), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_24__15_), .QN(n5529) );
  DFFR_X2 regBoiz_regfile_reg_18__15_ ( .D(n3979), .CK(clk), .RN(n6861), .Q(
        regBoiz_regfile_18__15_), .QN(n5528) );
  DFFR_X2 regBoiz_regfile_reg_16__15_ ( .D(n3977), .CK(clk), .RN(n6864), .Q(
        regBoiz_regfile_16__15_), .QN(n5527) );
  DFFR_X2 regBoiz_regfile_reg_2__15_ ( .D(n3963), .CK(clk), .RN(n6845), .Q(
        regBoiz_regfile_2__15_), .QN(n5526) );
  DFFR_X2 regBoiz_regfile_reg_0__15_ ( .D(n3961), .CK(clk), .RN(n6873), .Q(
        regBoiz_regfile_0__15_), .QN(n5525) );
  DFFRS_X1 ifBoi_pcOut_reg_26_ ( .D(n4583), .CK(clk), .RN(n3413), .SN(n3412), 
        .Q(iaddr[26]), .QN(n5520) );
  DFFR_X2 aluBoi_aluReg_45__regBoi_curData_reg ( .D(n4779), .CK(clk), .RN(
        n6889), .Q(daddr[1]), .QN(n5510) );
  DFFR_X2 ifBoi_reglol_66__regBoi_curData_reg ( .D(n4702), .CK(clk), .RN(n6911), .Q(ifOut_66_), .QN(n5508) );
  DFFR_X2 ifBoi_reglol_68__regBoi_curData_reg ( .D(n4690), .CK(clk), .RN(n6878), .Q(ifOut_68_), .QN(n5507) );
  DFFR_X2 ifBoi_reglol_72__regBoi_curData_reg ( .D(n4670), .CK(clk), .RN(n6898), .Q(ifOut_72_), .QN(n5506) );
  DFFR_X2 aluBoi_aluReg_58__regBoi_curData_reg ( .D(n4739), .CK(clk), .RN(
        n6890), .Q(daddr[14]), .QN(n5498) );
  DFFR_X2 aluBoi_aluReg_55__regBoi_curData_reg ( .D(n4745), .CK(clk), .RN(
        n6885), .Q(daddr[11]), .QN(n5497) );
  DFFR_X2 aluBoi_aluReg_54__regBoi_curData_reg ( .D(n4726), .CK(clk), .RN(
        n6890), .Q(daddr[10]), .QN(n5496) );
  DFFR_X2 aluBoi_aluReg_53__regBoi_curData_reg ( .D(n4730), .CK(clk), .RN(
        n6885), .Q(daddr[9]), .QN(n5495) );
  DFFR_X2 ifBoi_reglol_51__regBoi_curData_reg ( .D(n13595), .CK(clk), .RN(
        n6876), .Q(ifInst[19]), .QN(n5494) );
  DFFR_X2 ifBoi_reglol_49__regBoi_curData_reg ( .D(n13593), .CK(clk), .RN(
        n6897), .Q(ifInst[17]), .QN(n5493) );
  DFFR_X2 aluBoi_aluReg_56__regBoi_curData_reg ( .D(n4743), .CK(clk), .RN(
        n6890), .Q(daddr[12]), .QN(n5491) );
  DFFR_X2 ifBoi_reglol_70__regBoi_curData_reg ( .D(n4680), .CK(clk), .RN(n6898), .Q(ifOut_70_), .QN(n5490) );
  DFFR_X2 ifBoi_reglol_74__regBoi_curData_reg ( .D(n4662), .CK(clk), .RN(n6899), .Q(ifOut_74_), .QN(n5489) );
  DFFR_X2 aluBoi_aluReg_57__regBoi_curData_reg ( .D(n4741), .CK(clk), .RN(
        n6885), .Q(daddr[13]), .QN(n5488) );
  DFFR_X2 aluBoi_aluReg_52__regBoi_curData_reg ( .D(n4734), .CK(clk), .RN(
        n6889), .Q(daddr[8]), .QN(n5487) );
  DFFR_X2 ifBoi_reglol_47__regBoi_curData_reg ( .D(n13591), .CK(clk), .RN(
        n6897), .Q(ifInst[15]), .QN(n5485) );
  DFFR_X2 aluBoi_aluReg_59__regBoi_curData_reg ( .D(n4723), .CK(clk), .RN(
        n6885), .Q(daddr[15]), .QN(n5484) );
  DFFR_X2 ifBoi_reglol_41__regBoi_curData_reg ( .D(n13585), .CK(clk), .RN(
        n6897), .Q(ifInst[9]), .QN(n5481) );
  DFFR_X2 ifBoi_reglol_39__regBoi_curData_reg ( .D(n13583), .CK(clk), .RN(
        n6876), .Q(ifInst[7]), .QN(n5480) );
  DFFR_X2 ifBoi_reglol_50__regBoi_curData_reg ( .D(n13594), .CK(clk), .RN(
        n6897), .Q(ifInst[18]), .QN(n5479) );
  DFFR_X2 ifBoi_reglol_43__regBoi_curData_reg ( .D(n13587), .CK(clk), .RN(
        n6897), .Q(ifInst[11]), .QN(n5475) );
  DFFR_X2 ifBoi_reglol_45__regBoi_curData_reg ( .D(n13589), .CK(clk), .RN(
        n6897), .Q(ifInst[13]), .QN(n5473) );
  DFFR_X2 ifBoi_reglol_52__regBoi_curData_reg ( .D(n13596), .CK(clk), .RN(
        n6898), .Q(ifInst[20]), .QN(n5470) );
  DFFR_X2 ifBoi_reglol_40__regBoi_curData_reg ( .D(n13584), .CK(clk), .RN(
        n6876), .Q(ifInst[8]), .QN(n5469) );
  DFFR_X2 ifBoi_reglol_46__regBoi_curData_reg ( .D(n13590), .CK(clk), .RN(
        n6876), .Q(ifInst[14]), .QN(n5468) );
  DFFR_X2 ifBoi_reglol_48__regBoi_curData_reg ( .D(n13592), .CK(clk), .RN(
        n6876), .Q(ifInst[16]), .QN(n5467) );
  DFFR_X1 ifBoi_reglol_92__regBoi_curData_reg ( .D(n4572), .CK(clk), .RN(n6899), .Q(ifOut_92_), .QN(n5466) );
  DFFR_X2 ifBoi_reglol_42__regBoi_curData_reg ( .D(n13586), .CK(clk), .RN(
        n6876), .Q(ifInst[10]), .QN(n5465) );
  DFFR_X2 ifBoi_reglol_38__regBoi_curData_reg ( .D(n13582), .CK(clk), .RN(
        n6897), .Q(ifInst[6]), .QN(n5464) );
  DFFR_X2 ifBoi_reglol_44__regBoi_curData_reg ( .D(n13588), .CK(clk), .RN(
        n6876), .Q(ifInst[12]), .QN(n5463) );
  DFFR_X2 ifBoi_reglol_36__regBoi_curData_reg ( .D(n13580), .CK(clk), .RN(
        n6897), .Q(ifInst[4]), .QN(n5456) );
  DFFR_X2 ifBoi_reglol_62__regBoi_curData_reg ( .D(n13606), .CK(clk), .RN(
        n6905), .Q(ifInst[30]), .QN(n5455) );
  DFFR_X2 regBoiz_regfile_reg_19__21_ ( .D(n4178), .CK(clk), .RN(n6915), .Q(
        regBoiz_regfile_19__21_), .QN(n5402) );
  DFFR_X2 regBoiz_regfile_reg_26__14_ ( .D(n3954), .CK(clk), .RN(n6925), .Q(
        regBoiz_regfile_26__14_), .QN(n5401) );
  DFFR_X2 regBoiz_regfile_reg_18__14_ ( .D(n3946), .CK(clk), .RN(n6913), .Q(
        regBoiz_regfile_18__14_), .QN(n5400) );
  DFFR_X2 regBoiz_regfile_reg_10__14_ ( .D(n3938), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__14_), .QN(n5399) );
  DFFR_X2 regBoiz_regfile_reg_2__14_ ( .D(n3930), .CK(clk), .RN(n6931), .Q(
        regBoiz_regfile_2__14_), .QN(n5398) );
  DFFR_X2 regBoiz_regfile_reg_26__21_ ( .D(n4185), .CK(clk), .RN(n6926), .Q(
        regBoiz_regfile_26__21_), .QN(n5397) );
  DFFR_X2 regBoiz_regfile_reg_24__21_ ( .D(n4183), .CK(clk), .RN(n6923), .Q(
        regBoiz_regfile_24__21_), .QN(n5396) );
  DFFR_X2 idBoi_reggal_78__regBoi_curData_reg ( .D(n13615), .CK(clk), .RN(
        n6895), .Q(regBoiz_N17), .QN(n5389) );
  DFFR_X2 ifBoi_reglol_37__regBoi_curData_reg ( .D(n13581), .CK(clk), .RN(
        n6876), .Q(ifInst[5]), .QN(n5346) );
  DFFR_X2 idBoi_reggal_80__regBoi_curData_reg ( .D(n13617), .CK(clk), .RN(
        n6879), .QN(n5344) );
  DFFR_X2 ifBoi_reglol_35__regBoi_curData_reg ( .D(n13579), .CK(clk), .RN(
        n6877), .Q(ifInst[3]), .QN(n5343) );
  DFFR_X2 idBoi_reggal_77__regBoi_curData_reg ( .D(n13614), .CK(clk), .RN(
        n6879), .Q(regBoiz_N16), .QN(n5331) );
  DFFR_X2 aluBoi_aluReg_63__regBoi_curData_reg ( .D(n4746), .CK(clk), .RN(
        n6890), .Q(daddr[19]), .QN(n5323) );
  DFFR_X2 aluBoi_aluReg_60__regBoi_curData_reg ( .D(n4752), .CK(clk), .RN(
        n6884), .Q(daddr[16]), .QN(n5322) );
  DFFR_X2 idBoi_reggal_29__regBoi_curData_reg ( .D(n4791), .CK(clk), .RN(n6942), .Q(idOut_29_), .QN(n5314) );
  DFFR_X2 aluBoi_aluReg_41__regBoi_curData_reg ( .D(n4800), .CK(clk), .RN(
        n6889), .Q(aluRw[2]) );
  DFFR_X2 regBoiz_regfile_reg_14__27_ ( .D(n4371), .CK(clk), .RN(n6909), .Q(
        regBoiz_regfile_14__27_) );
  DFFR_X2 regBoiz_regfile_reg_30__20_ ( .D(n4156), .CK(clk), .RN(n6843), .Q(
        regBoiz_regfile_30__20_) );
  DFFR_X2 regBoiz_regfile_reg_23__8_ ( .D(n3753), .CK(clk), .RN(n6852), .Q(
        regBoiz_regfile_23__8_) );
  DFFR_X2 regBoiz_regfile_reg_10__27_ ( .D(n4367), .CK(clk), .RN(n6903), .Q(
        regBoiz_regfile_10__27_) );
  DFF_X1 aluBoi_multBoi_runProd_reg_54_ ( .D(aluBoi_multBoi_N60), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[50]) );
  DFFR_X2 aluBoi_aluReg_73__regBoi_curData_reg ( .D(n4773), .CK(clk), .RN(
        n6884), .Q(daddr[29]), .QN(n5327) );
  DFFR_X2 ifBoi_reglol_65__regBoi_curData_reg ( .D(n4707), .CK(clk), .RN(n6898), .Q(ifOut_65_) );
  DFF_X1 aluBoi_multBoi_runProd_reg_63_ ( .D(aluBoi_multBoi_N69), .CK(clk), 
        .Q(aluBoi_multBoi_temppp[59]) );
  INV_X4 U5099 ( .A(didMult), .ZN(net100619) );
  NAND2_X1 U5100 ( .A1(n8586), .A2(n6541), .ZN(n9072) );
  XNOR2_X1 U5101 ( .A(n8587), .B(n6541), .ZN(n9105) );
  INV_X2 U5102 ( .A(n6541), .ZN(n9635) );
  NAND2_X4 U5103 ( .A1(n6225), .A2(n6226), .ZN(n11126) );
  NAND2_X2 U5104 ( .A1(n11097), .A2(net361437), .ZN(n6225) );
  NOR3_X2 U5105 ( .A1(n11195), .A2(n11194), .A3(n11231), .ZN(n11198) );
  NOR2_X2 U5106 ( .A1(n11231), .A2(n11185), .ZN(n11061) );
  AOI21_X1 U5107 ( .B1(net360618), .B2(net360617), .A(net360619), .ZN(
        net360611) );
  OAI21_X2 U5108 ( .B1(net360611), .B2(n11678), .A(n11677), .ZN(net360604) );
  BUF_X16 U5109 ( .A(n12042), .Z(n4977) );
  INV_X2 U5110 ( .A(net361629), .ZN(n5783) );
  NOR2_X1 U5111 ( .A1(net361535), .A2(net361536), .ZN(n5777) );
  INV_X2 U5112 ( .A(net376076), .ZN(n4978) );
  INV_X1 U5113 ( .A(n12170), .ZN(n4979) );
  INV_X4 U5114 ( .A(n11425), .ZN(n11401) );
  XNOR2_X1 U5115 ( .A(n12427), .B(n12426), .ZN(n12432) );
  OAI21_X4 U5116 ( .B1(net359651), .B2(net359652), .A(net377513), .ZN(
        net359650) );
  INV_X2 U5117 ( .A(net359451), .ZN(net377513) );
  OAI21_X2 U5118 ( .B1(n7677), .B2(n7676), .A(n7675), .ZN(n4980) );
  NAND2_X2 U5119 ( .A1(n10951), .A2(n10950), .ZN(n4981) );
  OAI21_X2 U5120 ( .B1(n13706), .B2(n5947), .A(net368519), .ZN(n10951) );
  INV_X1 U5121 ( .A(n12301), .ZN(n4982) );
  INV_X2 U5122 ( .A(n4982), .ZN(n4983) );
  XNOR2_X1 U5123 ( .A(n6536), .B(n8762), .ZN(n9463) );
  NAND2_X1 U5124 ( .A1(n5288), .A2(n6536), .ZN(n9665) );
  NAND2_X1 U5125 ( .A1(net368215), .A2(n6536), .ZN(n10932) );
  INV_X2 U5126 ( .A(n9463), .ZN(n9468) );
  NAND2_X4 U5127 ( .A1(net376916), .A2(n6148), .ZN(n4984) );
  INV_X4 U5128 ( .A(n12088), .ZN(n4985) );
  INV_X8 U5129 ( .A(n12100), .ZN(n12088) );
  INV_X4 U5130 ( .A(n5982), .ZN(n6428) );
  OAI22_X2 U5131 ( .A1(n10189), .A2(net368447), .B1(n5033), .B2(net368187), 
        .ZN(n11440) );
  OAI21_X2 U5132 ( .B1(n5033), .B2(net368179), .A(n11451), .ZN(n11687) );
  XNOR2_X2 U5133 ( .A(n11612), .B(net377607), .ZN(n4987) );
  INV_X8 U5134 ( .A(n11777), .ZN(n11815) );
  AND2_X2 U5135 ( .A1(n11452), .A2(n11687), .ZN(n4988) );
  NAND2_X1 U5136 ( .A1(n11616), .A2(n11615), .ZN(n11617) );
  NAND4_X2 U5137 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n5266), .ZN(
        n12440) );
  INV_X1 U5138 ( .A(n11786), .ZN(n11802) );
  NAND2_X2 U5139 ( .A1(net360007), .A2(net360008), .ZN(net359524) );
  AND4_X2 U5140 ( .A1(net360273), .A2(n5483), .A3(net359533), .A4(net359535), 
        .ZN(n5342) );
  NAND3_X2 U5141 ( .A1(n11856), .A2(n11855), .A3(n11854), .ZN(n11859) );
  OAI211_X4 U5142 ( .C1(n12246), .C2(n12245), .A(n12243), .B(n12244), .ZN(
        n12393) );
  NAND2_X2 U5143 ( .A1(n11573), .A2(n11572), .ZN(n11575) );
  INV_X1 U5144 ( .A(n7526), .ZN(n4989) );
  INV_X2 U5145 ( .A(n4989), .ZN(n4990) );
  INV_X32 U5146 ( .A(n6251), .ZN(n10570) );
  INV_X1 U5147 ( .A(n12187), .ZN(n4991) );
  INV_X4 U5148 ( .A(n12252), .ZN(n12187) );
  XNOR2_X1 U5149 ( .A(n12172), .B(n12162), .ZN(n12068) );
  INV_X2 U5150 ( .A(n12174), .ZN(n12178) );
  BUF_X16 U5151 ( .A(n12047), .Z(n4994) );
  BUF_X32 U5152 ( .A(n12020), .Z(n4992) );
  XNOR2_X2 U5153 ( .A(n10883), .B(n10884), .ZN(n4993) );
  NAND2_X2 U5154 ( .A1(n10563), .A2(n10562), .ZN(n5892) );
  INV_X8 U5155 ( .A(n10927), .ZN(n10988) );
  INV_X8 U5156 ( .A(n7574), .ZN(n9829) );
  XNOR2_X2 U5157 ( .A(n4995), .B(net366989), .ZN(n6994) );
  NAND4_X1 U5158 ( .A1(n11340), .A2(net361053), .A3(n11367), .A4(n11341), .ZN(
        n4996) );
  XNOR2_X2 U5159 ( .A(n11336), .B(n11337), .ZN(n11341) );
  XNOR2_X2 U5160 ( .A(n10745), .B(n10827), .ZN(n4997) );
  OAI22_X4 U5161 ( .A1(n11731), .A2(net368467), .B1(net368211), .B2(n11833), 
        .ZN(n4998) );
  INV_X1 U5162 ( .A(n6061), .ZN(n11014) );
  NAND4_X2 U5163 ( .A1(n11179), .A2(n11181), .A3(n10892), .A4(n6536), .ZN(
        n4999) );
  NAND4_X2 U5164 ( .A1(n11179), .A2(n11181), .A3(n10892), .A4(n6536), .ZN(
        n10903) );
  NOR2_X2 U5165 ( .A1(n11388), .A2(n11387), .ZN(n11396) );
  NAND2_X2 U5166 ( .A1(n5948), .A2(n11478), .ZN(n5031) );
  INV_X2 U5167 ( .A(net369208), .ZN(n5242) );
  INV_X4 U5168 ( .A(n11949), .ZN(n6048) );
  NAND2_X2 U5169 ( .A1(n11933), .A2(net360299), .ZN(n12122) );
  INV_X2 U5170 ( .A(n12093), .ZN(n11922) );
  NOR2_X2 U5171 ( .A1(n6000), .A2(n11742), .ZN(n11743) );
  NAND3_X2 U5172 ( .A1(n11773), .A2(n11978), .A3(n11977), .ZN(n5000) );
  NAND3_X1 U5173 ( .A1(n11773), .A2(n11978), .A3(n11977), .ZN(n5001) );
  INV_X16 U5174 ( .A(n11772), .ZN(n11978) );
  NAND2_X4 U5175 ( .A1(n10479), .A2(n10478), .ZN(n5002) );
  OAI21_X2 U5176 ( .B1(n11653), .B2(n11652), .A(n11714), .ZN(n11753) );
  INV_X8 U5177 ( .A(n10836), .ZN(n5003) );
  INV_X4 U5178 ( .A(n10836), .ZN(n10971) );
  XNOR2_X2 U5179 ( .A(n12239), .B(n12081), .ZN(n5004) );
  INV_X4 U5180 ( .A(n5004), .ZN(n12282) );
  INV_X2 U5181 ( .A(n12081), .ZN(n12238) );
  INV_X8 U5182 ( .A(n10848), .ZN(n5005) );
  INV_X4 U5183 ( .A(n10848), .ZN(n10969) );
  XNOR2_X2 U5184 ( .A(n11864), .B(n5995), .ZN(n5006) );
  NAND2_X4 U5185 ( .A1(n5907), .A2(n10703), .ZN(n5007) );
  NAND2_X2 U5186 ( .A1(n11500), .A2(n11441), .ZN(n11407) );
  INV_X2 U5187 ( .A(n11483), .ZN(n6062) );
  XNOR2_X1 U5188 ( .A(n11483), .B(n6523), .ZN(n11546) );
  OAI21_X2 U5189 ( .B1(n11483), .B2(n6523), .A(n6521), .ZN(n11531) );
  NAND2_X2 U5190 ( .A1(net362257), .A2(net360821), .ZN(n10468) );
  NOR2_X2 U5191 ( .A1(n11626), .A2(n11388), .ZN(n5008) );
  INV_X4 U5192 ( .A(n12277), .ZN(n12371) );
  INV_X32 U5193 ( .A(net375310), .ZN(net378321) );
  XOR2_X2 U5194 ( .A(n12403), .B(n6212), .Z(n5009) );
  INV_X4 U5195 ( .A(n12402), .ZN(n6212) );
  AOI21_X2 U5196 ( .B1(n7790), .B2(n7789), .A(net366951), .ZN(n7794) );
  INV_X8 U5197 ( .A(n4984), .ZN(net359679) );
  OAI21_X2 U5198 ( .B1(n7828), .B2(n7827), .A(net366999), .ZN(n7829) );
  NAND2_X2 U5199 ( .A1(n4980), .A2(n9894), .ZN(n11183) );
  OAI22_X4 U5200 ( .A1(n11776), .A2(net368462), .B1(net368195), .B2(n11833), 
        .ZN(n11780) );
  AOI21_X4 U5201 ( .B1(n12530), .B2(n12531), .A(n12529), .ZN(n12533) );
  INV_X8 U5202 ( .A(n9790), .ZN(n10906) );
  NAND2_X1 U5203 ( .A1(ifOut_65_), .A2(idBoi_temPC_1_), .ZN(n9907) );
  NAND2_X1 U5204 ( .A1(ifOut_65_), .A2(n6582), .ZN(n12906) );
  OAI21_X2 U5205 ( .B1(n10396), .B2(n10397), .A(n9907), .ZN(n10385) );
  INV_X1 U5206 ( .A(n10280), .ZN(n5011) );
  INV_X4 U5207 ( .A(n5011), .ZN(n5012) );
  INV_X8 U5208 ( .A(n5459), .ZN(ifInst[0]) );
  OAI22_X1 U5209 ( .A1(n6602), .A2(n13459), .B1(n6597), .B2(n5459), .ZN(n13576) );
  INV_X1 U5210 ( .A(n10255), .ZN(n5014) );
  INV_X4 U5211 ( .A(n5014), .ZN(n5015) );
  INV_X8 U5212 ( .A(n5312), .ZN(ifInst[2]) );
  XOR2_X2 U5213 ( .A(n5508), .B(idBoi_temPC_2_), .Z(n10384) );
  NAND2_X1 U5214 ( .A1(n6581), .A2(ifInst[2]), .ZN(n13405) );
  OAI22_X1 U5215 ( .A1(n6602), .A2(n13461), .B1(n6594), .B2(n5312), .ZN(n13578) );
  XOR2_X1 U5216 ( .A(n10397), .B(n10396), .Z(n10398) );
  XNOR2_X1 U5217 ( .A(n10337), .B(n10336), .ZN(n10341) );
  XNOR2_X1 U5218 ( .A(n10308), .B(n10307), .ZN(n10311) );
  XNOR2_X1 U5219 ( .A(n5012), .B(n10279), .ZN(n10282) );
  XNOR2_X1 U5220 ( .A(n5015), .B(n10254), .ZN(n10257) );
  AOI222_X1 U5221 ( .A1(n12982), .A2(n13091), .B1(aluBoi_multBoi_temppp[16]), 
        .B2(net368069), .C1(n5316), .C2(aluBoi_imm32w_3_), .ZN(n13096) );
  INV_X4 U5222 ( .A(n11170), .ZN(aluBoi_multBoi_N50) );
  NOR2_X4 U5223 ( .A1(n9977), .A2(n9976), .ZN(n5017) );
  NOR2_X2 U5224 ( .A1(n9977), .A2(n9976), .ZN(n10045) );
  OAI221_X4 U5225 ( .B1(n9760), .B2(n9759), .C1(n9758), .C2(n13222), .A(n9757), 
        .ZN(n13182) );
  XNOR2_X2 U5226 ( .A(n10668), .B(n10671), .ZN(n10669) );
  XNOR2_X2 U5227 ( .A(n10671), .B(n5913), .ZN(n12317) );
  NAND2_X4 U5228 ( .A1(n10657), .A2(n10649), .ZN(n10671) );
  INV_X4 U5229 ( .A(net361309), .ZN(net359557) );
  NOR2_X2 U5230 ( .A1(n12223), .A2(net367631), .ZN(aluBoi_multBoi_N51) );
  NAND2_X4 U5231 ( .A1(n12498), .A2(net361306), .ZN(n10880) );
  NOR3_X2 U5232 ( .A1(net359552), .A2(net359553), .A3(net368481), .ZN(
        aluBoi_multBoi_N48) );
  OAI211_X1 U5233 ( .C1(net359557), .C2(n12499), .A(n12498), .B(net100619), 
        .ZN(n12500) );
  NAND2_X4 U5234 ( .A1(n12499), .A2(net359557), .ZN(n12498) );
  NAND2_X4 U5235 ( .A1(n10757), .A2(n5026), .ZN(n10859) );
  OAI21_X4 U5236 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n13238) );
  AOI222_X1 U5237 ( .A1(aluBoi_multBoi_temppp[25]), .A2(net368069), .B1(
        daddr[28]), .B2(n6609), .C1(n5316), .C2(aluBoi_imm32w_12_), .ZN(n13193) );
  INV_X4 U5238 ( .A(n10416), .ZN(n9610) );
  AOI22_X1 U5239 ( .A1(n9612), .A2(n10416), .B1(aluBoi_aluBoi_shft_srlout[6]), 
        .B2(n5381), .ZN(n9613) );
  INV_X1 U5240 ( .A(n8696), .ZN(n8662) );
  INV_X2 U5241 ( .A(n8882), .ZN(n5018) );
  BUF_X32 U5242 ( .A(n13269), .Z(n5019) );
  INV_X1 U5243 ( .A(n13255), .ZN(n13258) );
  NAND2_X4 U5244 ( .A1(n8706), .A2(n8705), .ZN(n8707) );
  AOI22_X1 U5245 ( .A1(n9633), .A2(n10415), .B1(aluBoi_aluBoi_shft_srlout[7]), 
        .B2(n5381), .ZN(n9634) );
  INV_X2 U5246 ( .A(n8587), .ZN(n8586) );
  INV_X8 U5247 ( .A(n6035), .ZN(n8701) );
  INV_X2 U5248 ( .A(n9492), .ZN(n5020) );
  XOR2_X2 U5249 ( .A(n6565), .B(n9492), .Z(n5021) );
  INV_X16 U5250 ( .A(n9677), .ZN(n6565) );
  INV_X8 U5251 ( .A(n10412), .ZN(n9492) );
  CLKBUF_X3 U5252 ( .A(n11937), .Z(n6015) );
  XNOR2_X2 U5253 ( .A(n6015), .B(aluBoi_multBoi_temppp[51]), .ZN(n5022) );
  NOR2_X2 U5254 ( .A1(n12333), .A2(net368481), .ZN(aluBoi_multBoi_N61) );
  MUX2_X1 U5255 ( .A(n8312), .B(n8311), .S(n6808), .Z(n8313) );
  AOI222_X1 U5256 ( .A1(aluBoi_multBoi_temppp[27]), .A2(net368069), .B1(
        daddr[30]), .B2(n6609), .C1(n5316), .C2(aluBoi_imm32w_14_), .ZN(n13230) );
  NOR3_X2 U5257 ( .A1(n5579), .A2(n13229), .A3(n13228), .ZN(n13232) );
  OAI21_X2 U5258 ( .B1(n13232), .B2(n13231), .A(n13230), .ZN(n4771) );
  BUF_X4 U5259 ( .A(net375910), .Z(net377824) );
  NOR2_X1 U5260 ( .A1(n5796), .A2(net377824), .ZN(net359521) );
  XNOR2_X2 U5261 ( .A(n6015), .B(aluBoi_multBoi_temppp[51]), .ZN(n5023) );
  INV_X4 U5262 ( .A(n5023), .ZN(net359540) );
  NOR2_X2 U5263 ( .A1(net359772), .A2(net359515), .ZN(net359904) );
  INV_X4 U5264 ( .A(n8883), .ZN(n8933) );
  NAND3_X2 U5265 ( .A1(n12509), .A2(net377689), .A3(net359537), .ZN(n12514) );
  INV_X32 U5266 ( .A(net369140), .ZN(net369147) );
  BUF_X4 U5267 ( .A(net369138), .Z(net369140) );
  AOI22_X1 U5268 ( .A1(n9494), .A2(n5020), .B1(aluBoi_aluBoi_shft_srlout[5]), 
        .B2(n5381), .ZN(n9495) );
  OAI21_X2 U5269 ( .B1(net359504), .B2(n12525), .A(net100619), .ZN(n12526) );
  NAND2_X2 U5270 ( .A1(net359680), .A2(n11971), .ZN(n11972) );
  NOR2_X2 U5271 ( .A1(n12335), .A2(n12334), .ZN(n12341) );
  NAND2_X4 U5272 ( .A1(n8724), .A2(n8723), .ZN(n9065) );
  XNOR2_X2 U5273 ( .A(n9756), .B(n9755), .ZN(n9758) );
  NAND4_X2 U5274 ( .A1(n12122), .A2(n11960), .A3(n12123), .A4(n11961), .ZN(
        n11962) );
  INV_X4 U5275 ( .A(n9199), .ZN(n6079) );
  OAI22_X4 U5276 ( .A1(n5305), .A2(n9117), .B1(n9116), .B2(n9115), .ZN(n9199)
         );
  INV_X8 U5277 ( .A(net359784), .ZN(net361266) );
  CLKBUF_X2 U5278 ( .A(net359492), .Z(net377979) );
  NOR2_X2 U5279 ( .A1(n12341), .A2(n12340), .ZN(aluBoi_multBoi_N65) );
  INV_X4 U5280 ( .A(net360284), .ZN(net360607) );
  NAND2_X2 U5281 ( .A1(n12505), .A2(n12506), .ZN(n5025) );
  NOR3_X2 U5282 ( .A1(net360278), .A2(n5801), .A3(net360279), .ZN(n5797) );
  NAND2_X2 U5283 ( .A1(n12520), .A2(n12519), .ZN(n12523) );
  NOR2_X4 U5284 ( .A1(n12527), .A2(n12526), .ZN(aluBoi_multBoi_N64) );
  NAND2_X4 U5285 ( .A1(net360607), .A2(net360606), .ZN(n12510) );
  INV_X2 U5286 ( .A(net360285), .ZN(net360606) );
  OAI21_X4 U5287 ( .B1(n10469), .B2(net368209), .A(n6117), .ZN(n10488) );
  XNOR2_X2 U5288 ( .A(aluBoi_multBoi_temppp[48]), .B(n11674), .ZN(n11436) );
  INV_X8 U5289 ( .A(net327826), .ZN(n11725) );
  INV_X8 U5290 ( .A(net377607), .ZN(net360550) );
  INV_X2 U5291 ( .A(net361838), .ZN(n5026) );
  INV_X4 U5292 ( .A(net361814), .ZN(net361838) );
  XNOR2_X2 U5293 ( .A(n11161), .B(n11337), .ZN(n5942) );
  NAND2_X2 U5294 ( .A1(net360632), .A2(net360626), .ZN(net361261) );
  INV_X8 U5295 ( .A(n11766), .ZN(n11729) );
  NAND2_X2 U5296 ( .A1(n11719), .A2(n11720), .ZN(n11766) );
  CLKBUF_X3 U5297 ( .A(n12423), .Z(n5027) );
  INV_X8 U5298 ( .A(net359507), .ZN(net359504) );
  AOI21_X2 U5299 ( .B1(n10448), .B2(n10449), .A(n5310), .ZN(n10450) );
  INV_X2 U5300 ( .A(n5891), .ZN(n5215) );
  INV_X4 U5301 ( .A(n12463), .ZN(n12436) );
  NAND2_X4 U5302 ( .A1(n5222), .A2(n5221), .ZN(net359488) );
  NAND2_X4 U5303 ( .A1(n12510), .A2(net359533), .ZN(n12505) );
  XNOR2_X2 U5304 ( .A(n11930), .B(n6013), .ZN(n5028) );
  NAND2_X2 U5305 ( .A1(net377576), .A2(net362050), .ZN(n10623) );
  AOI21_X4 U5306 ( .B1(n11165), .B2(n5226), .A(net361302), .ZN(n5029) );
  AOI21_X2 U5307 ( .B1(n11165), .B2(n5226), .A(net361302), .ZN(net361299) );
  NAND2_X2 U5308 ( .A1(n11321), .A2(n11354), .ZN(n5226) );
  XNOR2_X2 U5309 ( .A(n5000), .B(n6515), .ZN(n5030) );
  INV_X4 U5310 ( .A(net369206), .ZN(n5245) );
  OAI21_X4 U5311 ( .B1(n7501), .B2(net368548), .A(n7500), .ZN(n13522) );
  INV_X4 U5312 ( .A(n12015), .ZN(n11793) );
  INV_X8 U5313 ( .A(n11476), .ZN(n11478) );
  MUX2_X2 U5314 ( .A(regBoiz_regfile_2__27_), .B(regBoiz_regfile_10__27_), .S(
        net368782), .Z(n5809) );
  NAND2_X2 U5315 ( .A1(net359489), .A2(net377602), .ZN(n5221) );
  OAI22_X4 U5316 ( .A1(n7573), .A2(n7572), .B1(n7571), .B2(n7570), .ZN(n7574)
         );
  NAND2_X1 U5317 ( .A1(n7670), .A2(net367045), .ZN(n7572) );
  XNOR2_X2 U5318 ( .A(n11250), .B(n13521), .ZN(n5033) );
  NAND2_X4 U5319 ( .A1(n11372), .A2(n5977), .ZN(n5034) );
  NAND2_X2 U5320 ( .A1(n11299), .A2(n6525), .ZN(n11378) );
  AND2_X2 U5321 ( .A1(aluBoi_aluBoi_shft_sllout[15]), .A2(n5315), .ZN(n5035)
         );
  AOI22_X4 U5322 ( .A1(n9755), .A2(n9756), .B1(n9414), .B2(n5309), .ZN(n9768)
         );
  AND2_X2 U5323 ( .A1(n12215), .A2(net100619), .ZN(n5036) );
  NAND3_X4 U5324 ( .A1(n10721), .A2(n10616), .A3(n11229), .ZN(n5881) );
  INV_X2 U5325 ( .A(n11533), .ZN(n11571) );
  XNOR2_X1 U5326 ( .A(n11638), .B(n11751), .ZN(n11533) );
  AND3_X2 U5327 ( .A1(net368201), .A2(n10994), .A3(n10999), .ZN(n5037) );
  INV_X32 U5328 ( .A(n6593), .ZN(n6592) );
  INV_X8 U5329 ( .A(n13506), .ZN(n6593) );
  INV_X32 U5330 ( .A(n6592), .ZN(n6598) );
  AND2_X2 U5331 ( .A1(n12916), .A2(n5285), .ZN(n5038) );
  INV_X16 U5332 ( .A(n6591), .ZN(n6588) );
  INV_X8 U5333 ( .A(n6591), .ZN(n6590) );
  NAND2_X4 U5334 ( .A1(n6607), .A2(n5285), .ZN(n13430) );
  INV_X8 U5335 ( .A(n13363), .ZN(n6580) );
  NAND2_X2 U5336 ( .A1(n9994), .A2(n5285), .ZN(n10332) );
  INV_X8 U5337 ( .A(n10332), .ZN(n10286) );
  OAI22_X4 U5338 ( .A1(n11982), .A2(net368467), .B1(net368211), .B2(n12204), 
        .ZN(n5966) );
  OAI22_X4 U5339 ( .A1(n11731), .A2(net368467), .B1(net368211), .B2(n11833), 
        .ZN(n5895) );
  NAND2_X4 U5340 ( .A1(n11717), .A2(n11716), .ZN(n11805) );
  AND2_X2 U5341 ( .A1(n11609), .A2(n11610), .ZN(n5039) );
  INV_X16 U5342 ( .A(n10846), .ZN(n10955) );
  INV_X8 U5343 ( .A(n11643), .ZN(n6422) );
  AND2_X2 U5344 ( .A1(n4993), .A2(n6029), .ZN(n5040) );
  NAND2_X4 U5345 ( .A1(n11398), .A2(n11400), .ZN(n11281) );
  NAND2_X2 U5346 ( .A1(net361802), .A2(n6003), .ZN(n10816) );
  NAND2_X4 U5347 ( .A1(n11092), .A2(n11093), .ZN(n11037) );
  INV_X1 U5348 ( .A(n12274), .ZN(n6386) );
  INV_X4 U5349 ( .A(n12270), .ZN(n12272) );
  XOR2_X2 U5350 ( .A(n12347), .B(n12474), .Z(n5041) );
  AND2_X2 U5351 ( .A1(n12074), .A2(n12435), .ZN(n5042) );
  NAND2_X4 U5352 ( .A1(n11848), .A2(n11847), .ZN(n11856) );
  INV_X8 U5353 ( .A(n11749), .ZN(n11841) );
  INV_X4 U5354 ( .A(net361890), .ZN(net378420) );
  AND2_X2 U5355 ( .A1(n11103), .A2(n6429), .ZN(n5043) );
  NOR2_X4 U5356 ( .A1(net361539), .A2(net378420), .ZN(net361828) );
  INV_X4 U5357 ( .A(net361325), .ZN(n5836) );
  NAND2_X4 U5358 ( .A1(n11685), .A2(n11684), .ZN(n11960) );
  INV_X8 U5359 ( .A(n11913), .ZN(n11917) );
  AND2_X2 U5360 ( .A1(n5004), .A2(n12408), .ZN(n5044) );
  NOR2_X4 U5361 ( .A1(n12288), .A2(n12287), .ZN(n12283) );
  INV_X8 U5362 ( .A(n12241), .ZN(n12236) );
  INV_X16 U5363 ( .A(n12373), .ZN(n6392) );
  XOR2_X1 U5364 ( .A(net360235), .B(n5483), .Z(n5045) );
  AND3_X4 U5365 ( .A1(net361814), .A2(n11143), .A3(n11147), .ZN(n5046) );
  AND2_X4 U5366 ( .A1(net361292), .A2(net361293), .ZN(n5047) );
  AND2_X2 U5367 ( .A1(net359520), .A2(net359486), .ZN(n5048) );
  NAND2_X4 U5368 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  NAND2_X2 U5369 ( .A1(net360651), .A2(net360620), .ZN(n11435) );
  INV_X8 U5370 ( .A(net360996), .ZN(net360915) );
  AND2_X2 U5371 ( .A1(n12329), .A2(net100619), .ZN(n5049) );
  INV_X8 U5372 ( .A(n11301), .ZN(n11229) );
  NAND2_X2 U5373 ( .A1(net360904), .A2(net362257), .ZN(n10545) );
  INV_X4 U5374 ( .A(n5997), .ZN(n5050) );
  NAND2_X4 U5375 ( .A1(n5039), .A2(n11611), .ZN(n11612) );
  NAND2_X4 U5376 ( .A1(n5051), .A2(n5052), .ZN(n5053) );
  NAND2_X4 U5377 ( .A1(n11805), .A2(n5053), .ZN(n11636) );
  INV_X2 U5378 ( .A(n11717), .ZN(n5051) );
  INV_X4 U5379 ( .A(n11716), .ZN(n5052) );
  INV_X4 U5380 ( .A(n11796), .ZN(n5997) );
  NOR2_X4 U5381 ( .A1(n6420), .A2(n11608), .ZN(n11610) );
  NOR4_X2 U5382 ( .A1(n11625), .A2(n11624), .A3(n11636), .A4(n6553), .ZN(
        n11653) );
  INV_X8 U5383 ( .A(n11636), .ZN(n11796) );
  INV_X2 U5384 ( .A(n9791), .ZN(n7929) );
  AOI21_X4 U5385 ( .B1(n7920), .B2(n7919), .A(net366925), .ZN(n7921) );
  NAND2_X2 U5386 ( .A1(n7230), .A2(n7229), .ZN(n9801) );
  NAND2_X4 U5387 ( .A1(regBoiz_regfile_25__25_), .A2(n6787), .ZN(n7913) );
  NAND2_X2 U5388 ( .A1(net360904), .A2(net368498), .ZN(n10466) );
  NOR3_X4 U5389 ( .A1(net364898), .A2(net364899), .A3(net367041), .ZN(n5846)
         );
  NAND2_X2 U5390 ( .A1(n10711), .A2(n10710), .ZN(n5057) );
  NAND2_X4 U5391 ( .A1(n5055), .A2(n5056), .ZN(n5058) );
  NAND2_X4 U5392 ( .A1(n5057), .A2(n5058), .ZN(n10712) );
  INV_X8 U5393 ( .A(n10711), .ZN(n5055) );
  INV_X8 U5394 ( .A(n10710), .ZN(n5056) );
  NAND2_X1 U5395 ( .A1(n10708), .A2(net368201), .ZN(n10711) );
  NAND2_X2 U5396 ( .A1(net362224), .A2(n5843), .ZN(n5059) );
  NAND3_X1 U5397 ( .A1(net377695), .A2(n5839), .A3(n5060), .ZN(n5840) );
  INV_X2 U5398 ( .A(n5059), .ZN(n5060) );
  INV_X8 U5399 ( .A(n11594), .ZN(n11464) );
  OAI211_X4 U5400 ( .C1(n10575), .C2(net362172), .A(n10574), .B(net368215), 
        .ZN(n10576) );
  NAND2_X4 U5401 ( .A1(net362061), .A2(net362062), .ZN(n10622) );
  NAND2_X1 U5402 ( .A1(regBoiz_regfile_6__29_), .A2(n6770), .ZN(n181) );
  MUX2_X1 U5403 ( .A(regBoiz_regfile_6__29_), .B(regBoiz_regfile_7__29_), .S(
        net369157), .Z(n8264) );
  NAND2_X4 U5404 ( .A1(n6787), .A2(n8169), .ZN(n8170) );
  NAND4_X4 U5405 ( .A1(n5264), .A2(n5869), .A3(n10780), .A4(n11181), .ZN(
        n10815) );
  NAND2_X2 U5406 ( .A1(n7967), .A2(n5061), .ZN(n5062) );
  NAND2_X2 U5407 ( .A1(n7966), .A2(net366973), .ZN(n5063) );
  NAND2_X2 U5408 ( .A1(n5062), .A2(n5063), .ZN(net365100) );
  INV_X1 U5409 ( .A(net366973), .ZN(n5061) );
  INV_X4 U5410 ( .A(n6140), .ZN(n7966) );
  INV_X4 U5411 ( .A(n9786), .ZN(n9787) );
  NAND2_X4 U5412 ( .A1(n7968), .A2(net365099), .ZN(n9786) );
  NAND2_X2 U5413 ( .A1(n7226), .A2(n5064), .ZN(n5065) );
  NAND2_X1 U5414 ( .A1(n7225), .A2(net378321), .ZN(n5066) );
  NAND2_X2 U5415 ( .A1(n5065), .A2(n5066), .ZN(n7227) );
  INV_X1 U5416 ( .A(net378321), .ZN(n5064) );
  XNOR2_X2 U5417 ( .A(n10762), .B(n5102), .ZN(n10753) );
  INV_X8 U5418 ( .A(net375310), .ZN(net366935) );
  INV_X2 U5419 ( .A(net360254), .ZN(net360253) );
  NAND2_X4 U5420 ( .A1(n12359), .A2(n12358), .ZN(n12466) );
  NAND2_X4 U5421 ( .A1(regBoiz_regfile_27__25_), .A2(n6788), .ZN(n7919) );
  OAI21_X2 U5422 ( .B1(n7922), .B2(n7921), .A(net366969), .ZN(n7923) );
  INV_X16 U5423 ( .A(n13524), .ZN(n6542) );
  MUX2_X1 U5424 ( .A(regBoiz_regfile_14__20_), .B(regBoiz_regfile_30__20_), 
        .S(n6370), .Z(n7658) );
  INV_X8 U5425 ( .A(n11188), .ZN(n11298) );
  MUX2_X1 U5426 ( .A(n7224), .B(n7223), .S(net366981), .Z(n7225) );
  MUX2_X1 U5427 ( .A(regBoiz_regfile_14__8_), .B(regBoiz_regfile_15__8_), .S(
        net368800), .Z(n7223) );
  NAND2_X2 U5428 ( .A1(n7246), .A2(n7245), .ZN(n9799) );
  OAI21_X4 U5429 ( .B1(n5033), .B2(net368209), .A(n11284), .ZN(n11372) );
  INV_X8 U5430 ( .A(n6532), .ZN(n6533) );
  NAND4_X4 U5431 ( .A1(n6080), .A2(n10799), .A3(n10798), .A4(n10797), .ZN(
        n11144) );
  NAND2_X2 U5432 ( .A1(n7579), .A2(n8025), .ZN(n5234) );
  XNOR2_X1 U5433 ( .A(n11079), .B(n11204), .ZN(n11172) );
  INV_X4 U5434 ( .A(n11078), .ZN(n11077) );
  NAND2_X4 U5435 ( .A1(n11078), .A2(n11402), .ZN(n11206) );
  NAND2_X4 U5436 ( .A1(n7959), .A2(n9846), .ZN(n7960) );
  NAND2_X2 U5437 ( .A1(net359788), .A2(net361266), .ZN(net361262) );
  NAND2_X4 U5438 ( .A1(n7521), .A2(net367031), .ZN(n11056) );
  INV_X1 U5439 ( .A(net361830), .ZN(net378422) );
  AND2_X2 U5440 ( .A1(n12419), .A2(n12418), .ZN(n5068) );
  NAND2_X1 U5441 ( .A1(regBoiz_regfile_3__20_), .A2(n5069), .ZN(n5070) );
  NAND2_X1 U5442 ( .A1(regBoiz_regfile_19__20_), .A2(n6785), .ZN(n5071) );
  NAND2_X2 U5443 ( .A1(n5070), .A2(n5071), .ZN(n7655) );
  INV_X1 U5444 ( .A(n6785), .ZN(n5069) );
  NOR2_X2 U5445 ( .A1(n11551), .A2(n6553), .ZN(n11554) );
  NAND2_X1 U5446 ( .A1(n12205), .A2(net359942), .ZN(n5074) );
  NAND2_X4 U5447 ( .A1(n5072), .A2(n5073), .ZN(n5075) );
  NAND2_X2 U5448 ( .A1(n5074), .A2(n5075), .ZN(n12206) );
  INV_X4 U5449 ( .A(n12205), .ZN(n5072) );
  INV_X4 U5450 ( .A(net359942), .ZN(n5073) );
  NAND2_X1 U5451 ( .A1(net361902), .A2(n6040), .ZN(n5078) );
  NAND2_X4 U5452 ( .A1(n5076), .A2(n5077), .ZN(n5079) );
  NAND2_X4 U5453 ( .A1(n5078), .A2(n5079), .ZN(n11022) );
  INV_X2 U5454 ( .A(net361902), .ZN(n5076) );
  INV_X1 U5455 ( .A(n6040), .ZN(n5077) );
  NAND3_X2 U5456 ( .A1(n12031), .A2(n12123), .A3(n11566), .ZN(n5080) );
  INV_X4 U5457 ( .A(net377452), .ZN(net359942) );
  NOR2_X4 U5458 ( .A1(n12206), .A2(net367631), .ZN(aluBoi_multBoi_N66) );
  NAND2_X2 U5459 ( .A1(n8068), .A2(n5081), .ZN(n5082) );
  NAND2_X1 U5460 ( .A1(n8067), .A2(net366987), .ZN(n5083) );
  NAND2_X2 U5461 ( .A1(n5082), .A2(n5083), .ZN(n8069) );
  INV_X1 U5462 ( .A(net366987), .ZN(n5081) );
  NAND2_X2 U5463 ( .A1(n11797), .A2(n11798), .ZN(n11828) );
  XNOR2_X2 U5464 ( .A(net361537), .B(n5778), .ZN(n5776) );
  INV_X8 U5465 ( .A(n5944), .ZN(net365335) );
  NAND2_X1 U5466 ( .A1(regBoiz_regfile_18__22_), .A2(n5084), .ZN(n5085) );
  NAND2_X1 U5467 ( .A1(regBoiz_regfile_26__22_), .A2(n5242), .ZN(n5086) );
  NAND2_X2 U5468 ( .A1(n5085), .A2(n5086), .ZN(n7756) );
  INV_X1 U5469 ( .A(net375510), .ZN(n5084) );
  INV_X4 U5470 ( .A(n11254), .ZN(n11199) );
  NAND3_X1 U5471 ( .A1(net361491), .A2(n9829), .A3(n9830), .ZN(n9840) );
  INV_X8 U5472 ( .A(n11834), .ZN(n6154) );
  INV_X4 U5473 ( .A(n11806), .ZN(n6215) );
  INV_X8 U5474 ( .A(net360265), .ZN(n5804) );
  NAND4_X4 U5475 ( .A1(n5813), .A2(net377443), .A3(net361398), .A4(net361404), 
        .ZN(net361410) );
  INV_X4 U5476 ( .A(n12419), .ZN(n12420) );
  NAND2_X2 U5477 ( .A1(n9789), .A2(n10682), .ZN(n9790) );
  NOR2_X4 U5478 ( .A1(net359486), .A2(net359487), .ZN(n12529) );
  NAND2_X4 U5479 ( .A1(net360605), .A2(n6122), .ZN(n11665) );
  INV_X8 U5480 ( .A(n10596), .ZN(n10597) );
  NAND2_X4 U5481 ( .A1(n10595), .A2(n10594), .ZN(n10649) );
  INV_X8 U5482 ( .A(net375510), .ZN(net375867) );
  NAND2_X1 U5483 ( .A1(regBoiz_regfile_11__18_), .A2(n5087), .ZN(n5088) );
  NAND2_X1 U5484 ( .A1(regBoiz_regfile_27__18_), .A2(n6786), .ZN(n5089) );
  NAND2_X2 U5485 ( .A1(n5088), .A2(n5089), .ZN(n7586) );
  INV_X1 U5486 ( .A(n6786), .ZN(n5087) );
  NAND2_X2 U5487 ( .A1(n7998), .A2(n5090), .ZN(n5091) );
  NAND2_X1 U5488 ( .A1(n7997), .A2(net366987), .ZN(n5092) );
  NAND2_X2 U5489 ( .A1(n5091), .A2(n5092), .ZN(n7999) );
  INV_X1 U5490 ( .A(net366987), .ZN(n5090) );
  NAND2_X2 U5491 ( .A1(n7999), .A2(n9867), .ZN(net365033) );
  CLKBUF_X3 U5492 ( .A(n6783), .Z(n5093) );
  AND2_X4 U5493 ( .A1(n5094), .A2(n11182), .ZN(n11236) );
  AND3_X2 U5494 ( .A1(n11181), .A2(n11180), .A3(n11179), .ZN(n5094) );
  INV_X4 U5495 ( .A(n10564), .ZN(n5256) );
  NAND2_X1 U5496 ( .A1(regBoiz_regfile_14__27_), .A2(n6695), .ZN(n955) );
  MUX2_X1 U5497 ( .A(regBoiz_regfile_14__27_), .B(regBoiz_regfile_15__27_), 
        .S(net369161), .Z(n8197) );
  NAND3_X4 U5498 ( .A1(n6995), .A2(n6994), .A3(n6996), .ZN(n5944) );
  INV_X8 U5499 ( .A(n12134), .ZN(n12136) );
  INV_X1 U5500 ( .A(net377071), .ZN(net359766) );
  INV_X8 U5501 ( .A(n12336), .ZN(n12532) );
  NAND2_X2 U5502 ( .A1(n8041), .A2(n5095), .ZN(n5096) );
  NAND2_X1 U5503 ( .A1(n8040), .A2(net366977), .ZN(n5097) );
  NAND2_X2 U5504 ( .A1(n5096), .A2(n5097), .ZN(n8042) );
  INV_X1 U5505 ( .A(net366977), .ZN(n5095) );
  NAND2_X2 U5506 ( .A1(n8043), .A2(n8042), .ZN(n10478) );
  NAND2_X2 U5507 ( .A1(n7555), .A2(n5446), .ZN(n6110) );
  NAND2_X4 U5508 ( .A1(n10540), .A2(n10539), .ZN(net362159) );
  NOR2_X2 U5509 ( .A1(n11066), .A2(n10897), .ZN(n10898) );
  OAI21_X2 U5510 ( .B1(n11066), .B2(n10908), .A(n10973), .ZN(n10909) );
  NAND2_X2 U5511 ( .A1(n7242), .A2(n5098), .ZN(n5099) );
  NAND2_X1 U5512 ( .A1(n7241), .A2(net366939), .ZN(n5100) );
  NAND2_X2 U5513 ( .A1(n5099), .A2(n5100), .ZN(n7243) );
  INV_X1 U5514 ( .A(net366939), .ZN(n5098) );
  INV_X1 U5515 ( .A(net359494), .ZN(n5101) );
  INV_X1 U5516 ( .A(n6080), .ZN(n5102) );
  NAND2_X2 U5517 ( .A1(n7995), .A2(n5103), .ZN(n5104) );
  NAND2_X1 U5518 ( .A1(n7994), .A2(net366977), .ZN(n5105) );
  NAND2_X2 U5519 ( .A1(n5104), .A2(n5105), .ZN(n7996) );
  INV_X1 U5520 ( .A(net366977), .ZN(n5103) );
  NAND2_X2 U5521 ( .A1(n7996), .A2(n9846), .ZN(net365032) );
  INV_X4 U5522 ( .A(n12564), .ZN(n12566) );
  NAND2_X4 U5523 ( .A1(n10720), .A2(n10719), .ZN(n10828) );
  INV_X4 U5524 ( .A(n6783), .ZN(n5106) );
  INV_X4 U5525 ( .A(n5106), .ZN(n5107) );
  NAND2_X1 U5526 ( .A1(n10703), .A2(n9879), .ZN(n5108) );
  NAND2_X2 U5527 ( .A1(n5109), .A2(n6174), .ZN(n5936) );
  INV_X4 U5528 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U5529 ( .A1(n12009), .A2(n12105), .ZN(n5112) );
  NAND2_X2 U5530 ( .A1(n5110), .A2(n5111), .ZN(n5113) );
  NAND2_X4 U5531 ( .A1(n5112), .A2(n5113), .ZN(n12242) );
  INV_X2 U5532 ( .A(n12009), .ZN(n5110) );
  INV_X1 U5533 ( .A(n12105), .ZN(n5111) );
  NAND2_X2 U5534 ( .A1(n12285), .A2(n5134), .ZN(n12286) );
  BUF_X4 U5535 ( .A(n12127), .Z(n6034) );
  NAND2_X2 U5536 ( .A1(n5876), .A2(n6168), .ZN(n6170) );
  NAND2_X4 U5537 ( .A1(net367005), .A2(n7934), .ZN(n7938) );
  NAND2_X1 U5538 ( .A1(regBoiz_regfile_22__28_), .A2(n6727), .ZN(n654) );
  NAND2_X2 U5539 ( .A1(n5794), .A2(aluBoi_multBoi_temppp[49]), .ZN(n5116) );
  NAND2_X4 U5540 ( .A1(n5114), .A2(n5115), .ZN(n5117) );
  NAND2_X4 U5541 ( .A1(n5116), .A2(n5117), .ZN(net359913) );
  INV_X4 U5542 ( .A(n5794), .ZN(n5114) );
  INV_X4 U5543 ( .A(aluBoi_multBoi_temppp[49]), .ZN(n5115) );
  CLKBUF_X2 U5544 ( .A(net359913), .Z(net377800) );
  MUX2_X1 U5545 ( .A(regBoiz_regfile_2__28_), .B(regBoiz_regfile_18__28_), .S(
        n6370), .Z(n8040) );
  NOR2_X1 U5546 ( .A1(n12450), .A2(n12385), .ZN(n12388) );
  MUX2_X1 U5547 ( .A(n7554), .B(n7553), .S(net366971), .Z(n7555) );
  INV_X16 U5548 ( .A(net375310), .ZN(net366939) );
  AND2_X4 U5549 ( .A1(n5233), .A2(n5234), .ZN(n7596) );
  NAND2_X2 U5550 ( .A1(n7599), .A2(n5118), .ZN(n5119) );
  NAND2_X2 U5551 ( .A1(n7598), .A2(net366971), .ZN(n5120) );
  NAND2_X2 U5552 ( .A1(n5119), .A2(n5120), .ZN(n7600) );
  INV_X1 U5553 ( .A(net366971), .ZN(n5118) );
  AOI21_X2 U5554 ( .B1(n5959), .B2(n7600), .A(net367041), .ZN(n7613) );
  CLKBUF_X3 U5555 ( .A(n11130), .Z(n5121) );
  NAND2_X1 U5556 ( .A1(n10632), .A2(n10633), .ZN(n6169) );
  INV_X2 U5557 ( .A(n10633), .ZN(n6168) );
  INV_X4 U5558 ( .A(n10612), .ZN(n6201) );
  INV_X4 U5559 ( .A(n9890), .ZN(n7865) );
  NAND2_X2 U5560 ( .A1(n11059), .A2(n11192), .ZN(n11185) );
  NAND4_X2 U5561 ( .A1(n10783), .A2(net361801), .A3(n11059), .A4(n11192), .ZN(
        n10785) );
  BUF_X4 U5562 ( .A(net360604), .Z(net377817) );
  NAND2_X4 U5563 ( .A1(n12245), .A2(n6033), .ZN(n5134) );
  OAI21_X4 U5564 ( .B1(n11241), .B2(n11240), .A(n11239), .ZN(n5977) );
  OAI21_X4 U5565 ( .B1(n7930), .B2(n5310), .A(n9792), .ZN(n13524) );
  NAND2_X4 U5566 ( .A1(net361416), .A2(net369287), .ZN(n5122) );
  INV_X4 U5567 ( .A(n11819), .ZN(n12041) );
  NAND4_X4 U5568 ( .A1(n7596), .A2(n7594), .A3(n7595), .A4(n7593), .ZN(n9830)
         );
  NAND3_X2 U5569 ( .A1(n11686), .A2(n11960), .A3(n11912), .ZN(n11695) );
  INV_X4 U5570 ( .A(n5820), .ZN(n5821) );
  NAND2_X4 U5571 ( .A1(n9791), .A2(n9792), .ZN(n9794) );
  NAND2_X2 U5572 ( .A1(n9792), .A2(net368548), .ZN(n9793) );
  INV_X4 U5573 ( .A(n5145), .ZN(n5123) );
  NAND2_X1 U5574 ( .A1(regBoiz_regfile_15__16_), .A2(n6699), .ZN(n933) );
  NAND2_X1 U5575 ( .A1(n5029), .A2(net376800), .ZN(n5860) );
  INV_X2 U5576 ( .A(net361299), .ZN(n5859) );
  NAND3_X4 U5577 ( .A1(n11528), .A2(n11609), .A3(n11527), .ZN(n11529) );
  AND2_X2 U5578 ( .A1(n10631), .A2(n10688), .ZN(n5876) );
  NAND2_X2 U5579 ( .A1(n12075), .A2(n12076), .ZN(n12154) );
  NAND3_X1 U5580 ( .A1(n10746), .A2(n10689), .A3(net368201), .ZN(n10692) );
  NAND2_X2 U5581 ( .A1(n10746), .A2(n11071), .ZN(n10752) );
  NAND3_X2 U5582 ( .A1(n6552), .A2(n11553), .A3(n11534), .ZN(n11541) );
  INV_X4 U5583 ( .A(n6539), .ZN(n5260) );
  NOR2_X2 U5584 ( .A1(net359681), .A2(net359905), .ZN(n5864) );
  AOI21_X1 U5585 ( .B1(regBoiz_regfile_10__19_), .B2(net366949), .A(n6783), 
        .ZN(n7625) );
  NAND2_X4 U5586 ( .A1(n6288), .A2(n6289), .ZN(n8177) );
  INV_X8 U5587 ( .A(net362120), .ZN(net362114) );
  NAND2_X2 U5588 ( .A1(net359679), .A2(net359772), .ZN(net377900) );
  INV_X4 U5589 ( .A(net359486), .ZN(net359772) );
  NAND2_X2 U5590 ( .A1(n5229), .A2(n5230), .ZN(net362135) );
  OAI21_X2 U5591 ( .B1(n10528), .B2(n5002), .A(n10526), .ZN(net362178) );
  NAND2_X2 U5592 ( .A1(n7283), .A2(n5124), .ZN(n5125) );
  NAND2_X1 U5593 ( .A1(n7282), .A2(net366927), .ZN(n5126) );
  NAND2_X2 U5594 ( .A1(n5125), .A2(n5126), .ZN(n7291) );
  INV_X1 U5595 ( .A(net366927), .ZN(n5124) );
  NOR2_X4 U5596 ( .A1(n5816), .A2(net359497), .ZN(net377784) );
  NAND2_X1 U5597 ( .A1(n12156), .A2(n12358), .ZN(n5129) );
  NAND2_X2 U5598 ( .A1(n5127), .A2(n5128), .ZN(n5130) );
  NAND2_X4 U5599 ( .A1(n5129), .A2(n5130), .ZN(n12158) );
  INV_X4 U5600 ( .A(n12156), .ZN(n5127) );
  INV_X1 U5601 ( .A(n12358), .ZN(n5128) );
  NAND2_X2 U5602 ( .A1(n5382), .A2(n5131), .ZN(n5132) );
  NAND2_X1 U5603 ( .A1(n5588), .A2(net376331), .ZN(n5133) );
  NAND2_X2 U5604 ( .A1(n5132), .A2(n5133), .ZN(n7955) );
  INV_X1 U5605 ( .A(net376331), .ZN(n5131) );
  OAI21_X1 U5606 ( .B1(net361000), .B2(net361001), .A(net361002), .ZN(n5788)
         );
  NAND2_X4 U5607 ( .A1(n11158), .A2(net378368), .ZN(net361007) );
  INV_X4 U5608 ( .A(net361013), .ZN(net378368) );
  NAND2_X2 U5609 ( .A1(n10761), .A2(n10800), .ZN(n6135) );
  NAND2_X4 U5610 ( .A1(n10914), .A2(n5151), .ZN(n11194) );
  INV_X2 U5611 ( .A(n10914), .ZN(n10916) );
  OAI21_X2 U5612 ( .B1(n5332), .B2(n11177), .A(n11176), .ZN(n11213) );
  INV_X8 U5613 ( .A(n11921), .ZN(n11923) );
  INV_X4 U5614 ( .A(n10823), .ZN(n6046) );
  INV_X1 U5615 ( .A(net376077), .ZN(n5135) );
  NAND2_X2 U5616 ( .A1(n11268), .A2(n11267), .ZN(n11269) );
  NAND3_X2 U5617 ( .A1(n11400), .A2(n5939), .A3(n11283), .ZN(n11267) );
  XNOR2_X1 U5618 ( .A(n10858), .B(n11154), .ZN(n11167) );
  INV_X4 U5619 ( .A(n11154), .ZN(n11157) );
  NOR2_X2 U5620 ( .A1(n11391), .A2(n5212), .ZN(n11392) );
  NOR2_X2 U5621 ( .A1(n6059), .A2(n6275), .ZN(n12124) );
  NAND3_X2 U5622 ( .A1(net361491), .A2(n9832), .A3(n9831), .ZN(n9839) );
  OAI211_X4 U5623 ( .C1(n11394), .C2(n11281), .A(n11393), .B(n11392), .ZN(
        n11395) );
  INV_X8 U5624 ( .A(n10702), .ZN(n10720) );
  INV_X8 U5625 ( .A(n11112), .ZN(n13706) );
  NAND2_X2 U5626 ( .A1(n10792), .A2(n13706), .ZN(n10793) );
  INV_X8 U5627 ( .A(n10446), .ZN(n8052) );
  NOR2_X4 U5628 ( .A1(n12543), .A2(net359418), .ZN(n12544) );
  INV_X16 U5629 ( .A(net345751), .ZN(net362287) );
  OAI21_X4 U5630 ( .B1(n10517), .B2(n10516), .A(n10515), .ZN(n10625) );
  OAI211_X2 U5631 ( .C1(net377462), .C2(net360926), .A(net361023), .B(n5792), 
        .ZN(net360919) );
  OAI21_X4 U5632 ( .B1(n6380), .B2(n10514), .A(n5902), .ZN(n10515) );
  INV_X2 U5633 ( .A(n11125), .ZN(n11098) );
  XNOR2_X2 U5634 ( .A(n12256), .B(n12348), .ZN(n12164) );
  NAND2_X4 U5635 ( .A1(net362238), .A2(net362237), .ZN(net377080) );
  OAI21_X4 U5636 ( .B1(net362269), .B2(net368548), .A(net362265), .ZN(
        net362238) );
  INV_X4 U5637 ( .A(net361404), .ZN(net361401) );
  AOI21_X4 U5638 ( .B1(n12276), .B2(n12357), .A(n12361), .ZN(n12277) );
  INV_X4 U5639 ( .A(n12069), .ZN(n12170) );
  INV_X4 U5640 ( .A(n9787), .ZN(n5872) );
  INV_X16 U5641 ( .A(n6539), .ZN(n10892) );
  NAND2_X2 U5642 ( .A1(n12143), .A2(n12142), .ZN(n5138) );
  NAND2_X4 U5643 ( .A1(n5136), .A2(n5137), .ZN(n5139) );
  NAND2_X4 U5644 ( .A1(n5138), .A2(n5139), .ZN(net359507) );
  INV_X8 U5645 ( .A(n12143), .ZN(n5136) );
  INV_X4 U5646 ( .A(n12142), .ZN(n5137) );
  NAND2_X2 U5647 ( .A1(net359507), .A2(n12144), .ZN(net359675) );
  INV_X2 U5648 ( .A(n5944), .ZN(n5140) );
  NOR2_X4 U5649 ( .A1(n11230), .A2(n10897), .ZN(n10899) );
  AOI22_X4 U5650 ( .A1(n7589), .A2(n7670), .B1(n7588), .B2(n5446), .ZN(n7594)
         );
  OAI21_X2 U5651 ( .B1(n12300), .B2(n12299), .A(n12298), .ZN(n12302) );
  NAND2_X1 U5652 ( .A1(n11435), .A2(n11678), .ZN(n5143) );
  NAND2_X4 U5653 ( .A1(n5141), .A2(n5142), .ZN(n5144) );
  NAND2_X4 U5654 ( .A1(n5143), .A2(n5144), .ZN(n11668) );
  INV_X4 U5655 ( .A(n11435), .ZN(n5141) );
  INV_X2 U5656 ( .A(n11678), .ZN(n5142) );
  NAND2_X4 U5657 ( .A1(n11108), .A2(n11107), .ZN(n11110) );
  XOR2_X2 U5658 ( .A(net360474), .B(n5894), .Z(n5920) );
  INV_X32 U5659 ( .A(net366905), .ZN(net376374) );
  INV_X4 U5660 ( .A(n9819), .ZN(n7521) );
  INV_X8 U5661 ( .A(net361831), .ZN(n5145) );
  INV_X4 U5662 ( .A(net361831), .ZN(net376139) );
  XOR2_X2 U5663 ( .A(n12580), .B(n12478), .Z(n5146) );
  XOR2_X2 U5664 ( .A(n12477), .B(n5146), .Z(n12479) );
  NAND2_X2 U5665 ( .A1(n12279), .A2(n12189), .ZN(n5149) );
  NAND2_X4 U5666 ( .A1(n5147), .A2(n5148), .ZN(n5150) );
  NAND2_X4 U5667 ( .A1(n5149), .A2(n5150), .ZN(n12360) );
  INV_X1 U5668 ( .A(n12279), .ZN(n5147) );
  INV_X4 U5669 ( .A(n12189), .ZN(n5148) );
  INV_X1 U5670 ( .A(n12583), .ZN(n12478) );
  AOI211_X4 U5671 ( .C1(n12198), .C2(n5888), .A(n12360), .B(n12197), .ZN(
        n12202) );
  INV_X8 U5672 ( .A(n12360), .ZN(n12361) );
  NAND2_X2 U5673 ( .A1(n10503), .A2(n10608), .ZN(n10507) );
  OAI21_X4 U5674 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(n5151) );
  NAND2_X1 U5675 ( .A1(n10745), .A2(n10827), .ZN(n5154) );
  NAND2_X4 U5676 ( .A1(n5152), .A2(n5153), .ZN(n5155) );
  NAND2_X4 U5677 ( .A1(n5154), .A2(n5155), .ZN(n10835) );
  INV_X2 U5678 ( .A(n10745), .ZN(n5152) );
  INV_X2 U5679 ( .A(n10827), .ZN(n5153) );
  INV_X4 U5680 ( .A(n10835), .ZN(n10717) );
  NAND2_X2 U5681 ( .A1(n7305), .A2(n5156), .ZN(n5157) );
  NAND2_X1 U5682 ( .A1(n7304), .A2(net376077), .ZN(n5158) );
  NAND2_X2 U5683 ( .A1(n5157), .A2(n5158), .ZN(n7306) );
  INV_X1 U5684 ( .A(net376077), .ZN(n5156) );
  INV_X8 U5685 ( .A(net376076), .ZN(net376077) );
  NAND2_X1 U5686 ( .A1(n7306), .A2(n5093), .ZN(n6328) );
  INV_X4 U5687 ( .A(net375618), .ZN(n5159) );
  INV_X8 U5688 ( .A(net376223), .ZN(net375618) );
  NAND2_X2 U5689 ( .A1(n7545), .A2(n5160), .ZN(n5161) );
  NAND2_X1 U5690 ( .A1(n7544), .A2(net366969), .ZN(n5162) );
  NAND2_X2 U5691 ( .A1(n5161), .A2(n5162), .ZN(n7546) );
  INV_X1 U5692 ( .A(net366969), .ZN(n5160) );
  AOI22_X2 U5693 ( .A1(n8039), .A2(n7547), .B1(n8025), .B2(n7546), .ZN(n7564)
         );
  INV_X1 U5694 ( .A(n13533), .ZN(n11067) );
  NAND3_X2 U5695 ( .A1(n10729), .A2(n11197), .A3(net368213), .ZN(n10731) );
  NAND2_X1 U5696 ( .A1(n7512), .A2(n5163), .ZN(n5164) );
  NAND2_X1 U5697 ( .A1(n7513), .A2(n5275), .ZN(n5165) );
  NAND2_X2 U5698 ( .A1(n5164), .A2(n5165), .ZN(n9818) );
  INV_X1 U5699 ( .A(n5275), .ZN(n5163) );
  INV_X4 U5700 ( .A(net378321), .ZN(n5275) );
  NAND2_X1 U5701 ( .A1(net360904), .A2(n13533), .ZN(n11176) );
  NAND2_X4 U5702 ( .A1(n10776), .A2(n10777), .ZN(n5166) );
  NAND2_X1 U5703 ( .A1(n10774), .A2(n10775), .ZN(n5169) );
  NAND2_X4 U5704 ( .A1(n5167), .A2(n5168), .ZN(n5170) );
  NAND2_X4 U5705 ( .A1(n5169), .A2(n5170), .ZN(n10776) );
  INV_X2 U5706 ( .A(n10774), .ZN(n5167) );
  INV_X4 U5707 ( .A(n10775), .ZN(n5168) );
  INV_X4 U5708 ( .A(net376574), .ZN(n5171) );
  INV_X8 U5709 ( .A(net369202), .ZN(net376574) );
  INV_X16 U5710 ( .A(net369210), .ZN(net369200) );
  NAND2_X1 U5711 ( .A1(n11868), .A2(n11867), .ZN(n11998) );
  INV_X8 U5712 ( .A(net362237), .ZN(net362233) );
  NAND3_X2 U5713 ( .A1(net362268), .A2(net362265), .A3(net377481), .ZN(n5819)
         );
  INV_X8 U5714 ( .A(net361670), .ZN(net361802) );
  INV_X8 U5715 ( .A(net366905), .ZN(net366885) );
  NAND2_X2 U5716 ( .A1(n11837), .A2(n11838), .ZN(n11844) );
  INV_X4 U5717 ( .A(n5826), .ZN(n5827) );
  NAND4_X2 U5718 ( .A1(net369286), .A2(n6071), .A3(n11129), .A4(n11130), .ZN(
        n11131) );
  INV_X8 U5719 ( .A(n10559), .ZN(n6245) );
  INV_X2 U5720 ( .A(n11581), .ZN(n5175) );
  NAND2_X4 U5721 ( .A1(n10781), .A2(n10782), .ZN(n11193) );
  INV_X4 U5722 ( .A(net375867), .ZN(net378494) );
  BUF_X8 U5723 ( .A(net360919), .Z(net377947) );
  NAND3_X2 U5724 ( .A1(n5135), .A2(n7830), .A3(n7829), .ZN(n7831) );
  OAI21_X1 U5725 ( .B1(n7822), .B2(n7821), .A(net366967), .ZN(n7830) );
  INV_X2 U5726 ( .A(n11629), .ZN(n11596) );
  NAND2_X2 U5727 ( .A1(n7744), .A2(n5172), .ZN(n5173) );
  NAND2_X1 U5728 ( .A1(n7743), .A2(net366973), .ZN(n5174) );
  NAND2_X2 U5729 ( .A1(n5173), .A2(n5174), .ZN(n9847) );
  INV_X1 U5730 ( .A(net366973), .ZN(n5172) );
  INV_X4 U5731 ( .A(n9847), .ZN(n7745) );
  OAI222_X2 U5732 ( .A1(n9852), .A2(n9851), .B1(n9850), .B2(n9849), .C1(n9848), 
        .C2(n9847), .ZN(n9874) );
  NAND2_X1 U5733 ( .A1(n11581), .A2(n11557), .ZN(n5177) );
  NAND2_X4 U5734 ( .A1(n5175), .A2(n5176), .ZN(n5178) );
  NAND2_X2 U5735 ( .A1(n5177), .A2(n5178), .ZN(n11559) );
  INV_X4 U5736 ( .A(n11557), .ZN(n5176) );
  INV_X1 U5737 ( .A(n11582), .ZN(n11557) );
  NAND2_X4 U5738 ( .A1(n12080), .A2(n12079), .ZN(n12155) );
  NOR2_X1 U5739 ( .A1(n5310), .A2(n6793), .ZN(n7246) );
  NAND2_X2 U5740 ( .A1(n12045), .A2(n12044), .ZN(n12050) );
  MUX2_X1 U5741 ( .A(regBoiz_regfile_18__16_), .B(regBoiz_regfile_26__16_), 
        .S(net368782), .Z(n7508) );
  INV_X16 U5742 ( .A(net368782), .ZN(net375929) );
  NAND2_X2 U5743 ( .A1(regBoiz_regfile_12__31_), .A2(net368782), .ZN(n6287) );
  INV_X32 U5744 ( .A(net366901), .ZN(net368782) );
  NAND2_X2 U5745 ( .A1(n8071), .A2(n5179), .ZN(n5180) );
  NAND2_X1 U5746 ( .A1(n8070), .A2(net366977), .ZN(n5181) );
  NAND2_X2 U5747 ( .A1(n5180), .A2(n5181), .ZN(n8072) );
  INV_X1 U5748 ( .A(net366977), .ZN(n5179) );
  NOR2_X2 U5749 ( .A1(n5182), .A2(n5183), .ZN(n5184) );
  NOR2_X2 U5750 ( .A1(n5184), .A2(n10443), .ZN(n10449) );
  INV_X4 U5751 ( .A(n10444), .ZN(n5182) );
  INV_X4 U5752 ( .A(n10445), .ZN(n5183) );
  NOR2_X1 U5753 ( .A1(net367041), .A2(n6782), .ZN(n10445) );
  INV_X4 U5754 ( .A(n10442), .ZN(n10443) );
  INV_X4 U5755 ( .A(n10976), .ZN(n10987) );
  INV_X1 U5756 ( .A(n11855), .ZN(n5185) );
  INV_X2 U5757 ( .A(n5185), .ZN(n5186) );
  OAI222_X4 U5758 ( .A1(n7940), .A2(n7970), .B1(n7939), .B2(n7938), .C1(n7937), 
        .C2(n7936), .ZN(n7954) );
  NAND2_X4 U5759 ( .A1(n11753), .A2(n11752), .ZN(n11847) );
  NAND3_X2 U5760 ( .A1(n9843), .A2(n9844), .A3(n9845), .ZN(n5187) );
  NAND2_X4 U5761 ( .A1(n5188), .A2(n9842), .ZN(n11721) );
  INV_X4 U5762 ( .A(n5187), .ZN(n5188) );
  INV_X8 U5763 ( .A(net367013), .ZN(net367007) );
  INV_X8 U5764 ( .A(net359916), .ZN(net376581) );
  AND3_X2 U5765 ( .A1(n11052), .A2(n6531), .A3(net361491), .ZN(n5443) );
  NAND2_X2 U5766 ( .A1(n8164), .A2(n5189), .ZN(n5190) );
  NAND2_X1 U5767 ( .A1(n8163), .A2(net366987), .ZN(n5191) );
  NAND2_X2 U5768 ( .A1(n5190), .A2(n5191), .ZN(n8171) );
  INV_X1 U5769 ( .A(net366987), .ZN(n5189) );
  BUF_X4 U5770 ( .A(n11992), .Z(n6419) );
  OAI22_X1 U5771 ( .A1(n6024), .A2(net375527), .B1(n6025), .B2(net366995), 
        .ZN(n6023) );
  NAND4_X4 U5772 ( .A1(n11040), .A2(n11038), .A3(n11039), .A4(net361372), .ZN(
        n11080) );
  XNOR2_X2 U5773 ( .A(n11432), .B(n11745), .ZN(n11434) );
  OAI22_X1 U5774 ( .A1(n12166), .A2(net368446), .B1(n6049), .B2(net368187), 
        .ZN(n12279) );
  INV_X2 U5775 ( .A(n12255), .ZN(n12348) );
  NAND2_X4 U5776 ( .A1(n11871), .A2(n11875), .ZN(n11756) );
  NOR2_X4 U5777 ( .A1(net368498), .A2(n10536), .ZN(n10537) );
  NAND2_X2 U5778 ( .A1(net361027), .A2(n5192), .ZN(n5193) );
  NAND2_X4 U5779 ( .A1(n5193), .A2(n5862), .ZN(net360926) );
  INV_X1 U5780 ( .A(net361028), .ZN(n5192) );
  NAND2_X1 U5781 ( .A1(n11432), .A2(n11318), .ZN(n5196) );
  NAND2_X4 U5782 ( .A1(n5194), .A2(n5195), .ZN(n5197) );
  NAND2_X4 U5783 ( .A1(n5196), .A2(n5197), .ZN(net361030) );
  INV_X2 U5784 ( .A(n11432), .ZN(n5194) );
  INV_X4 U5785 ( .A(n11318), .ZN(n5195) );
  XNOR2_X1 U5786 ( .A(n6064), .B(n11317), .ZN(n11318) );
  NAND2_X2 U5787 ( .A1(net361031), .A2(net361030), .ZN(net361029) );
  MUX2_X1 U5788 ( .A(regBoiz_regfile_19__27_), .B(regBoiz_regfile_27__27_), 
        .S(net376077), .Z(n7971) );
  INV_X2 U5789 ( .A(net360620), .ZN(net360619) );
  NAND2_X2 U5790 ( .A1(n11977), .A2(n5286), .ZN(n11980) );
  CLKBUF_X3 U5791 ( .A(n11976), .Z(n5286) );
  OAI221_X4 U5792 ( .B1(n12275), .B2(n12274), .C1(n12273), .C2(n12272), .A(
        n12358), .ZN(n12276) );
  INV_X4 U5793 ( .A(n11278), .ZN(n11394) );
  NAND2_X4 U5794 ( .A1(n5198), .A2(n5199), .ZN(n5200) );
  NAND2_X4 U5795 ( .A1(n5200), .A2(n11492), .ZN(n11861) );
  INV_X4 U5796 ( .A(n11493), .ZN(n5198) );
  INV_X4 U5797 ( .A(n11421), .ZN(n5199) );
  INV_X2 U5798 ( .A(n11491), .ZN(n11492) );
  INV_X8 U5799 ( .A(n5781), .ZN(n5782) );
  NAND2_X2 U5800 ( .A1(n12532), .A2(net359766), .ZN(net359762) );
  INV_X4 U5801 ( .A(n11464), .ZN(n5202) );
  NAND2_X2 U5802 ( .A1(n11595), .A2(n11594), .ZN(n11628) );
  INV_X2 U5803 ( .A(n11401), .ZN(n5203) );
  INV_X4 U5804 ( .A(n5203), .ZN(n5204) );
  NAND2_X2 U5805 ( .A1(n7378), .A2(n5205), .ZN(n5206) );
  NAND2_X1 U5806 ( .A1(n7377), .A2(n6785), .ZN(n5207) );
  NAND2_X2 U5807 ( .A1(n5206), .A2(n5207), .ZN(n7379) );
  INV_X1 U5808 ( .A(n6785), .ZN(n5205) );
  OAI22_X1 U5809 ( .A1(n7358), .A2(net375717), .B1(n7357), .B2(net367043), 
        .ZN(n7359) );
  AOI22_X2 U5810 ( .A1(regBoiz_regfile_13__12_), .A2(net367003), .B1(
        regBoiz_regfile_15__12_), .B2(net366985), .ZN(n7357) );
  INV_X1 U5811 ( .A(n5935), .ZN(n11223) );
  NAND2_X4 U5812 ( .A1(n6442), .A2(n10958), .ZN(n10952) );
  AND2_X2 U5813 ( .A1(net361491), .A2(n11053), .ZN(n5208) );
  AND2_X2 U5814 ( .A1(n5906), .A2(n5208), .ZN(n5921) );
  NAND2_X1 U5815 ( .A1(n7527), .A2(n5209), .ZN(n5210) );
  NAND2_X1 U5816 ( .A1(n4990), .A2(net378321), .ZN(n5211) );
  NAND2_X2 U5817 ( .A1(n5210), .A2(n5211), .ZN(n5906) );
  INV_X1 U5818 ( .A(net378321), .ZN(n5209) );
  NAND2_X2 U5819 ( .A1(n11053), .A2(n5906), .ZN(n7528) );
  INV_X4 U5820 ( .A(n11302), .ZN(n11247) );
  OAI22_X4 U5821 ( .A1(n11991), .A2(net368462), .B1(net368195), .B2(n12204), 
        .ZN(n12048) );
  INV_X8 U5822 ( .A(n6095), .ZN(n11640) );
  INV_X2 U5823 ( .A(n11474), .ZN(n5212) );
  NAND2_X2 U5824 ( .A1(n6183), .A2(n6184), .ZN(n5935) );
  NAND2_X1 U5825 ( .A1(n5204), .A2(n11377), .ZN(n5213) );
  NOR2_X4 U5826 ( .A1(n12170), .A2(n5214), .ZN(n12181) );
  INV_X8 U5827 ( .A(n5911), .ZN(n5214) );
  NAND2_X2 U5828 ( .A1(n5891), .A2(net377607), .ZN(n5217) );
  NAND2_X2 U5829 ( .A1(n5215), .A2(n5216), .ZN(n5218) );
  NAND2_X2 U5830 ( .A1(n5217), .A2(n5218), .ZN(n11881) );
  INV_X1 U5831 ( .A(net377607), .ZN(n5216) );
  INV_X4 U5832 ( .A(n12167), .ZN(n12171) );
  INV_X1 U5833 ( .A(net359470), .ZN(net359651) );
  XOR2_X1 U5834 ( .A(n11501), .B(n11702), .Z(n11704) );
  XNOR2_X1 U5835 ( .A(n11501), .B(n11702), .ZN(n11857) );
  NOR4_X2 U5836 ( .A1(n10930), .A2(n6093), .A3(net368211), .A4(n11249), .ZN(
        n10934) );
  NAND2_X4 U5837 ( .A1(n6198), .A2(n10928), .ZN(n10972) );
  NAND2_X4 U5838 ( .A1(n10820), .A2(n10819), .ZN(n10883) );
  NAND2_X4 U5839 ( .A1(n10884), .A2(n10883), .ZN(n11036) );
  NAND2_X4 U5840 ( .A1(n11396), .A2(n11395), .ZN(n11441) );
  INV_X1 U5841 ( .A(n5880), .ZN(n11896) );
  NAND2_X2 U5842 ( .A1(n11191), .A2(n9828), .ZN(n5945) );
  OAI221_X4 U5843 ( .B1(n11870), .B2(n6249), .C1(n11852), .C2(n11851), .A(
        n11871), .ZN(n11853) );
  NAND2_X4 U5844 ( .A1(n5219), .A2(n5220), .ZN(n5222) );
  INV_X4 U5845 ( .A(net359489), .ZN(n5219) );
  INV_X4 U5846 ( .A(net377602), .ZN(n5220) );
  XNOR2_X1 U5847 ( .A(net361268), .B(n5685), .ZN(n5223) );
  NOR2_X4 U5848 ( .A1(net359488), .A2(net368481), .ZN(aluBoi_multBoi_N68) );
  NOR2_X2 U5849 ( .A1(n11877), .A2(n11876), .ZN(n11878) );
  NAND2_X4 U5850 ( .A1(net377081), .A2(net362239), .ZN(n5842) );
  AOI21_X2 U5851 ( .B1(n11811), .B2(n11816), .A(n11810), .ZN(n11831) );
  AOI211_X4 U5852 ( .C1(n11804), .C2(n11803), .A(n11802), .B(n11801), .ZN(
        n11811) );
  NAND2_X1 U5853 ( .A1(n11531), .A2(n11530), .ZN(n11655) );
  NAND2_X4 U5854 ( .A1(net368215), .A2(n11199), .ZN(n11062) );
  OAI21_X4 U5855 ( .B1(n5823), .B2(net361270), .A(net361271), .ZN(net361268)
         );
  INV_X1 U5856 ( .A(net361324), .ZN(n5224) );
  INV_X2 U5857 ( .A(n5224), .ZN(n5225) );
  INV_X16 U5858 ( .A(net376223), .ZN(net367043) );
  MUX2_X1 U5859 ( .A(regBoiz_regfile_22__8_), .B(regBoiz_regfile_23__8_), .S(
        net376223), .Z(n7233) );
  MUX2_X1 U5860 ( .A(regBoiz_regfile_30__0_), .B(regBoiz_regfile_31__0_), .S(
        net376223), .Z(n6984) );
  NAND2_X1 U5861 ( .A1(net378103), .A2(net362140), .ZN(n5229) );
  NAND2_X2 U5862 ( .A1(n5227), .A2(n5228), .ZN(n5230) );
  INV_X4 U5863 ( .A(net378103), .ZN(n5227) );
  INV_X1 U5864 ( .A(net362140), .ZN(n5228) );
  INV_X2 U5865 ( .A(n8162), .ZN(n8163) );
  BUF_X4 U5866 ( .A(n10855), .Z(n5769) );
  INV_X4 U5867 ( .A(n11524), .ZN(n5231) );
  INV_X8 U5868 ( .A(n6519), .ZN(n11524) );
  INV_X32 U5869 ( .A(n6526), .ZN(n6527) );
  NAND2_X2 U5870 ( .A1(regBoiz_regfile_28__14_), .A2(net366939), .ZN(n7443) );
  NAND2_X4 U5871 ( .A1(n10996), .A2(n6067), .ZN(n10997) );
  INV_X4 U5872 ( .A(net361320), .ZN(net361302) );
  INV_X2 U5873 ( .A(n11630), .ZN(n5232) );
  INV_X8 U5874 ( .A(n13536), .ZN(n6540) );
  INV_X2 U5875 ( .A(n11824), .ZN(n11799) );
  NOR2_X1 U5876 ( .A1(n11796), .A2(n11824), .ZN(n11621) );
  NAND2_X2 U5877 ( .A1(n8039), .A2(n7580), .ZN(n5233) );
  NAND2_X2 U5878 ( .A1(n6047), .A2(n11495), .ZN(n11429) );
  NAND2_X1 U5879 ( .A1(n11313), .A2(n11312), .ZN(n11431) );
  INV_X2 U5880 ( .A(n6535), .ZN(n11003) );
  NAND2_X1 U5881 ( .A1(regBoiz_regfile_21__29_), .A2(n5235), .ZN(n5236) );
  NAND2_X1 U5882 ( .A1(regBoiz_regfile_29__29_), .A2(net377166), .ZN(n5237) );
  NAND2_X2 U5883 ( .A1(n5236), .A2(n5237), .ZN(n8062) );
  INV_X1 U5884 ( .A(net377166), .ZN(n5235) );
  NAND2_X2 U5885 ( .A1(n8062), .A2(n5238), .ZN(n5239) );
  NAND2_X1 U5886 ( .A1(n8061), .A2(net366987), .ZN(n5240) );
  NAND2_X2 U5887 ( .A1(n5239), .A2(n5240), .ZN(n8063) );
  INV_X1 U5888 ( .A(net366987), .ZN(n5238) );
  NAND2_X2 U5889 ( .A1(n8063), .A2(net366933), .ZN(n10438) );
  NAND2_X2 U5890 ( .A1(regBoiz_regfile_19__28_), .A2(n6370), .ZN(n6138) );
  NAND3_X1 U5891 ( .A1(net366907), .A2(net366919), .A3(net366965), .ZN(n8007)
         );
  NAND2_X2 U5892 ( .A1(net366933), .A2(net366907), .ZN(n8106) );
  CLKBUF_X3 U5893 ( .A(n10552), .Z(n6380) );
  INV_X4 U5894 ( .A(net362342), .ZN(net375876) );
  NAND2_X4 U5895 ( .A1(n8066), .A2(net366953), .ZN(n10439) );
  NAND2_X2 U5896 ( .A1(net359752), .A2(net377611), .ZN(n5811) );
  INV_X2 U5897 ( .A(net377611), .ZN(net362485) );
  INV_X1 U5898 ( .A(n10913), .ZN(n5241) );
  NAND2_X1 U5899 ( .A1(regBoiz_regfile_24__27_), .A2(net369202), .ZN(n5243) );
  NAND2_X2 U5900 ( .A1(regBoiz_regfile_16__27_), .A2(net369208), .ZN(n5244) );
  NAND2_X2 U5901 ( .A1(n5243), .A2(n5244), .ZN(n6371) );
  CLKBUF_X3 U5902 ( .A(n12359), .Z(n5888) );
  NAND3_X2 U5903 ( .A1(n12392), .A2(n12375), .A3(aluBoi_multBoi_temppp[59]), 
        .ZN(n12306) );
  INV_X8 U5904 ( .A(net361433), .ZN(net361416) );
  INV_X2 U5905 ( .A(n8157), .ZN(n5972) );
  NOR2_X2 U5906 ( .A1(n6000), .A2(n11494), .ZN(n11498) );
  INV_X1 U5907 ( .A(n11615), .ZN(n6060) );
  NAND2_X1 U5908 ( .A1(net362240), .A2(net361984), .ZN(n5841) );
  NOR2_X4 U5909 ( .A1(n11178), .A2(n11207), .ZN(n5246) );
  OAI21_X2 U5910 ( .B1(n6425), .B2(n11400), .A(n11283), .ZN(n11207) );
  NAND2_X4 U5911 ( .A1(n11912), .A2(n6098), .ZN(n11953) );
  NOR2_X4 U5912 ( .A1(n12463), .A2(n12191), .ZN(n12192) );
  INV_X16 U5913 ( .A(n11722), .ZN(n11305) );
  INV_X8 U5914 ( .A(net361358), .ZN(net361746) );
  NAND2_X4 U5915 ( .A1(n7896), .A2(net375506), .ZN(n9791) );
  OR2_X2 U5916 ( .A1(n5247), .A2(net376541), .ZN(n5280) );
  INV_X2 U5917 ( .A(net376076), .ZN(net375980) );
  INV_X16 U5918 ( .A(net376374), .ZN(net376541) );
  NAND2_X4 U5919 ( .A1(n6195), .A2(n11330), .ZN(n6197) );
  NAND2_X2 U5920 ( .A1(n11347), .A2(n11346), .ZN(n6196) );
  OR2_X2 U5921 ( .A1(n6194), .A2(n10791), .ZN(n5889) );
  NAND2_X1 U5922 ( .A1(regBoiz_regfile_18__28_), .A2(n6709), .ZN(n820) );
  INV_X2 U5923 ( .A(n10527), .ZN(n10508) );
  NAND2_X4 U5924 ( .A1(n7879), .A2(n7878), .ZN(n7895) );
  NOR2_X2 U5925 ( .A1(n10912), .A2(n10913), .ZN(n10921) );
  INV_X4 U5926 ( .A(net359501), .ZN(net359499) );
  XNOR2_X2 U5927 ( .A(net360513), .B(n6215), .ZN(n11732) );
  NOR2_X4 U5928 ( .A1(n10519), .A2(n6115), .ZN(n10525) );
  INV_X16 U5929 ( .A(net376417), .ZN(n5248) );
  INV_X32 U5930 ( .A(net368781), .ZN(net376417) );
  NAND2_X4 U5931 ( .A1(n6135), .A2(n6136), .ZN(n10763) );
  MUX2_X2 U5932 ( .A(n5930), .B(n7955), .S(n5249), .Z(n7956) );
  INV_X32 U5933 ( .A(net366973), .ZN(n5249) );
  NAND2_X4 U5934 ( .A1(n7514), .A2(net375506), .ZN(n11055) );
  INV_X4 U5935 ( .A(n5900), .ZN(n7514) );
  NAND2_X4 U5936 ( .A1(n5250), .A2(n5251), .ZN(n5252) );
  NAND2_X2 U5937 ( .A1(n11613), .A2(n5252), .ZN(n11708) );
  INV_X4 U5938 ( .A(n11463), .ZN(n5250) );
  INV_X4 U5939 ( .A(n11462), .ZN(n5251) );
  INV_X8 U5940 ( .A(n11708), .ZN(n6552) );
  NOR2_X4 U5941 ( .A1(n6251), .A2(net368195), .ZN(n5253) );
  NOR2_X4 U5942 ( .A1(n10561), .A2(n5254), .ZN(n10565) );
  INV_X4 U5943 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U5944 ( .A1(n10564), .A2(n10565), .ZN(n5257) );
  NAND2_X4 U5945 ( .A1(n5255), .A2(n5256), .ZN(n5258) );
  NAND2_X4 U5946 ( .A1(n5257), .A2(n5258), .ZN(n5871) );
  INV_X2 U5947 ( .A(n10565), .ZN(n5255) );
  NOR2_X2 U5948 ( .A1(n5892), .A2(net375435), .ZN(n10564) );
  INV_X16 U5949 ( .A(n6529), .ZN(n11191) );
  NOR2_X4 U5950 ( .A1(net368462), .A2(n5260), .ZN(n5259) );
  INV_X4 U5951 ( .A(n5259), .ZN(n10924) );
  INV_X32 U5952 ( .A(net368462), .ZN(net360904) );
  NAND2_X4 U5953 ( .A1(n9846), .A2(n8177), .ZN(n8178) );
  NAND2_X1 U5954 ( .A1(regBoiz_regfile_8__28_), .A2(n5261), .ZN(n5262) );
  NAND2_X1 U5955 ( .A1(regBoiz_regfile_24__28_), .A2(n6783), .ZN(n5263) );
  NAND2_X2 U5956 ( .A1(n5262), .A2(n5263), .ZN(n8027) );
  INV_X1 U5957 ( .A(n6783), .ZN(n5261) );
  NAND3_X2 U5958 ( .A1(n5883), .A2(net362253), .A3(n10508), .ZN(n10509) );
  NAND2_X2 U5959 ( .A1(n10779), .A2(n10778), .ZN(n5264) );
  INV_X4 U5960 ( .A(n5883), .ZN(n5265) );
  INV_X8 U5961 ( .A(n10528), .ZN(n5883) );
  NAND2_X4 U5962 ( .A1(n11048), .A2(n5442), .ZN(n11043) );
  OAI21_X1 U5963 ( .B1(net361512), .B2(n5882), .A(n10989), .ZN(n10954) );
  NAND2_X2 U5964 ( .A1(n11477), .A2(n11187), .ZN(n11607) );
  INV_X8 U5965 ( .A(n11800), .ZN(n11801) );
  NAND2_X2 U5966 ( .A1(n5283), .A2(n5284), .ZN(n12592) );
  NAND2_X4 U5967 ( .A1(n10623), .A2(n10622), .ZN(n10628) );
  NAND2_X1 U5968 ( .A1(n11366), .A2(n11367), .ZN(net361001) );
  NAND3_X4 U5969 ( .A1(n6244), .A2(n12017), .A3(n12013), .ZN(n5266) );
  NAND3_X2 U5970 ( .A1(n6244), .A2(n12017), .A3(n12013), .ZN(n12433) );
  NAND2_X2 U5971 ( .A1(n11278), .A2(n6029), .ZN(n11009) );
  NAND2_X1 U5972 ( .A1(n9879), .A2(n10703), .ZN(n5267) );
  NAND2_X2 U5973 ( .A1(n5268), .A2(n6174), .ZN(n10781) );
  INV_X4 U5974 ( .A(n5267), .ZN(n5268) );
  NAND2_X1 U5975 ( .A1(n11113), .A2(n11129), .ZN(n11039) );
  NAND2_X1 U5976 ( .A1(n12241), .A2(n12240), .ZN(n5270) );
  NAND2_X2 U5977 ( .A1(n12236), .A2(n5269), .ZN(n5271) );
  NAND2_X2 U5978 ( .A1(n5270), .A2(n5271), .ZN(n12386) );
  INV_X1 U5979 ( .A(n12240), .ZN(n5269) );
  OAI21_X2 U5980 ( .B1(net368181), .B2(n12204), .A(n12203), .ZN(n12240) );
  NAND2_X4 U5981 ( .A1(n11968), .A2(n11967), .ZN(n12148) );
  INV_X8 U5982 ( .A(n10707), .ZN(n10719) );
  OAI22_X4 U5983 ( .A1(n5007), .A2(n10706), .B1(n10705), .B2(n10770), .ZN(
        n10707) );
  NAND2_X4 U5984 ( .A1(n11030), .A2(n10856), .ZN(net361548) );
  INV_X1 U5985 ( .A(net361835), .ZN(net361830) );
  NAND3_X2 U5986 ( .A1(n6048), .A2(n5418), .A3(n11963), .ZN(n11965) );
  AND2_X4 U5987 ( .A1(n11945), .A2(n11944), .ZN(n5418) );
  NOR2_X4 U5988 ( .A1(net359487), .A2(net359486), .ZN(n5272) );
  INV_X2 U5989 ( .A(n11019), .ZN(n6006) );
  NAND2_X4 U5990 ( .A1(n11836), .A2(n11931), .ZN(n11963) );
  INV_X4 U5991 ( .A(n11901), .ZN(n11931) );
  INV_X16 U5992 ( .A(n10726), .ZN(n10722) );
  INV_X4 U5993 ( .A(n11010), .ZN(n11008) );
  NAND2_X4 U5994 ( .A1(n10993), .A2(n10992), .ZN(n11085) );
  NAND3_X2 U5995 ( .A1(n11046), .A2(n10991), .A3(n10941), .ZN(n11010) );
  INV_X8 U5996 ( .A(n12290), .ZN(n12291) );
  INV_X8 U5997 ( .A(net368903), .ZN(net376642) );
  INV_X8 U5998 ( .A(net376642), .ZN(net376063) );
  INV_X4 U5999 ( .A(n11137), .ZN(n11135) );
  NAND2_X4 U6000 ( .A1(n11047), .A2(n11046), .ZN(n11050) );
  NOR2_X4 U6001 ( .A1(n11741), .A2(n11740), .ZN(n11744) );
  NOR3_X4 U6002 ( .A1(n11963), .A2(n11952), .A3(n11951), .ZN(n11948) );
  BUF_X4 U6003 ( .A(n11036), .Z(n5882) );
  NAND3_X2 U6004 ( .A1(n10961), .A2(n6029), .A3(n11035), .ZN(n10963) );
  NAND2_X1 U6005 ( .A1(n10703), .A2(net368548), .ZN(n9887) );
  MUX2_X2 U6006 ( .A(n7505), .B(n7504), .S(net366969), .Z(n7506) );
  INV_X2 U6007 ( .A(n6106), .ZN(n5274) );
  INV_X8 U6008 ( .A(net360282), .ZN(net360007) );
  INV_X8 U6009 ( .A(n10521), .ZN(n10510) );
  INV_X8 U6010 ( .A(n12237), .ZN(n12401) );
  INV_X4 U6011 ( .A(net361357), .ZN(net361748) );
  NAND2_X1 U6012 ( .A1(n10435), .A2(n5275), .ZN(n5276) );
  NAND2_X1 U6013 ( .A1(n10434), .A2(net378321), .ZN(n5277) );
  NAND2_X2 U6014 ( .A1(n5276), .A2(n5277), .ZN(n10444) );
  NAND2_X1 U6015 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  BUF_X4 U6016 ( .A(net360605), .Z(net377791) );
  OAI21_X4 U6017 ( .B1(n10510), .B2(net377937), .A(net362297), .ZN(n10683) );
  INV_X1 U6018 ( .A(net361532), .ZN(net361885) );
  BUF_X8 U6019 ( .A(net361056), .Z(net377550) );
  NAND3_X4 U6020 ( .A1(n10540), .A2(n10487), .A3(n10539), .ZN(net362327) );
  INV_X8 U6021 ( .A(n11867), .ZN(n11876) );
  INV_X8 U6022 ( .A(net368787), .ZN(net375510) );
  NOR2_X4 U6023 ( .A1(n11949), .A2(n11946), .ZN(n11888) );
  AND2_X2 U6024 ( .A1(n11550), .A2(n5008), .ZN(n6108) );
  INV_X4 U6025 ( .A(n10815), .ZN(n10783) );
  XNOR2_X2 U6026 ( .A(n11086), .B(n11085), .ZN(n11087) );
  NAND2_X1 U6027 ( .A1(regBoiz_regfile_6__16_), .A2(n5278), .ZN(n5279) );
  NAND2_X2 U6028 ( .A1(n5279), .A2(n5280), .ZN(n7504) );
  INV_X4 U6029 ( .A(net375980), .ZN(n5278) );
  NAND2_X1 U6030 ( .A1(n12591), .A2(n12590), .ZN(n5283) );
  NAND2_X4 U6031 ( .A1(n5281), .A2(n5282), .ZN(n5284) );
  INV_X4 U6032 ( .A(n12591), .ZN(n5281) );
  INV_X4 U6033 ( .A(n12590), .ZN(n5282) );
  NOR2_X4 U6034 ( .A1(n12592), .A2(net368481), .ZN(aluBoi_multBoi_N70) );
  NOR2_X4 U6035 ( .A1(n11301), .A2(n5945), .ZN(n11307) );
  BUF_X32 U6036 ( .A(n13303), .Z(n5285) );
  INV_X8 U6037 ( .A(didKill), .ZN(n13303) );
  INV_X4 U6038 ( .A(n9904), .ZN(n5287) );
  INV_X2 U6039 ( .A(n9904), .ZN(n9940) );
  NAND2_X1 U6040 ( .A1(n6575), .A2(aluBoi_aluBoi_shft_sraout[31]), .ZN(n9996)
         );
  NAND2_X1 U6041 ( .A1(aluBoi_aluBoi_shft_sraout[31]), .A2(n12944), .ZN(n13510) );
  OAI21_X1 U6042 ( .B1(n6562), .B2(n9723), .A(aluBoi_aluBoi_shft_sraout[31]), 
        .ZN(n9726) );
  OAI21_X1 U6043 ( .B1(aluBoi_aluBoi_shft_sraout[31]), .B2(n6564), .A(n6561), 
        .ZN(n9724) );
  NAND2_X1 U6044 ( .A1(net359603), .A2(aluBoi_aluBoi_shft_sraout[31]), .ZN(
        n12458) );
  NAND2_X1 U6045 ( .A1(net359752), .A2(aluBoi_aluBoi_shft_sraout[31]), .ZN(
        n12343) );
  INV_X2 U6046 ( .A(aluBoi_aluBoi_shft_sraout[31]), .ZN(n12251) );
  INV_X2 U6047 ( .A(aluBoi_aluBoi_shft_sraout[31]), .ZN(n12184) );
  INV_X16 U6048 ( .A(aluBoi_aluBoi_shft_sraout[31]), .ZN(n12183) );
  NAND2_X1 U6049 ( .A1(regBoiz_regfile_7__6_), .A2(n6772), .ZN(n139) );
  NAND2_X2 U6050 ( .A1(n6493), .A2(n6494), .ZN(n7183) );
  MUX2_X1 U6051 ( .A(n7156), .B(n7155), .S(net366967), .Z(n7157) );
  NAND2_X2 U6052 ( .A1(n9798), .A2(n9797), .ZN(n9811) );
  MUX2_X1 U6053 ( .A(n7295), .B(n7294), .S(net366979), .Z(n7296) );
  INV_X16 U6054 ( .A(n5310), .ZN(net361491) );
  INV_X8 U6055 ( .A(n9899), .ZN(n11977) );
  INV_X8 U6056 ( .A(net368681), .ZN(net368786) );
  INV_X16 U6057 ( .A(net368786), .ZN(net368787) );
  NAND4_X4 U6058 ( .A1(n10844), .A2(n6435), .A3(n10958), .A4(net378405), .ZN(
        n10847) );
  NAND2_X4 U6059 ( .A1(n11958), .A2(n11957), .ZN(n11968) );
  INV_X2 U6060 ( .A(n11000), .ZN(n11001) );
  NOR3_X4 U6061 ( .A1(n11217), .A2(n11216), .A3(n11215), .ZN(n11228) );
  NOR2_X4 U6062 ( .A1(n11044), .A2(n5970), .ZN(n11047) );
  NOR3_X4 U6063 ( .A1(n11886), .A2(n11949), .A3(n11928), .ZN(n11887) );
  INV_X8 U6064 ( .A(n12112), .ZN(n11949) );
  INV_X2 U6065 ( .A(n12416), .ZN(n6436) );
  MUX2_X1 U6066 ( .A(regBoiz_regfile_7__16_), .B(regBoiz_regfile_15__16_), .S(
        net375510), .Z(n7524) );
  NAND3_X4 U6067 ( .A1(n11055), .A2(n11056), .A3(n6787), .ZN(n7529) );
  OAI22_X2 U6068 ( .A1(net378420), .A2(net361536), .B1(net361889), .B2(
        net378420), .ZN(n5806) );
  XNOR2_X2 U6069 ( .A(n12285), .B(n12144), .ZN(n12143) );
  OAI21_X4 U6070 ( .B1(n12130), .B2(n12141), .A(n12140), .ZN(n12131) );
  OAI21_X4 U6071 ( .B1(n12141), .B2(n12130), .A(n12140), .ZN(n12142) );
  NOR2_X4 U6072 ( .A1(n6041), .A2(n12292), .ZN(n11964) );
  XNOR2_X2 U6073 ( .A(n11680), .B(n11667), .ZN(n12508) );
  NAND3_X4 U6074 ( .A1(n5819), .A2(net362264), .A3(net360821), .ZN(net362237)
         );
  NAND2_X1 U6075 ( .A1(n10715), .A2(net361949), .ZN(n10716) );
  NAND2_X2 U6076 ( .A1(regBoiz_regfile_12__29_), .A2(net369204), .ZN(n6126) );
  INV_X16 U6077 ( .A(net369206), .ZN(net369204) );
  NAND2_X4 U6078 ( .A1(n11941), .A2(n11944), .ZN(n11930) );
  NAND2_X4 U6079 ( .A1(n11672), .A2(n11673), .ZN(net360285) );
  OAI22_X4 U6080 ( .A1(n11644), .A2(n11645), .B1(n11644), .B2(n6423), .ZN(
        n11650) );
  NAND2_X4 U6081 ( .A1(net360283), .A2(net375910), .ZN(net360282) );
  OAI221_X4 U6082 ( .B1(net360284), .B2(net360285), .C1(n5342), .C2(net360287), 
        .A(net360288), .ZN(net360283) );
  XNOR2_X1 U6083 ( .A(n12182), .B(n12183), .ZN(n12459) );
  NAND2_X1 U6084 ( .A1(n6608), .A2(n5285), .ZN(n13363) );
  NAND2_X1 U6085 ( .A1(regBoiz_regfile_23__6_), .A2(n6728), .ZN(n612) );
  NAND2_X1 U6086 ( .A1(regBoiz_regfile_27__6_), .A2(n6743), .ZN(n477) );
  MUX2_X2 U6087 ( .A(regBoiz_regfile_26__6_), .B(regBoiz_regfile_27__6_), .S(
        net375717), .Z(n7173) );
  INV_X16 U6088 ( .A(net366901), .ZN(net366899) );
  NAND2_X2 U6089 ( .A1(n13303), .A2(n12916), .ZN(difKill) );
  MUX2_X1 U6090 ( .A(n7118), .B(n7117), .S(net375650), .Z(n7119) );
  NAND2_X4 U6091 ( .A1(n7121), .A2(net361491), .ZN(n9797) );
  NAND2_X2 U6092 ( .A1(n9903), .A2(idOut_32_), .ZN(n6239) );
  NAND2_X4 U6093 ( .A1(n9901), .A2(n9902), .ZN(n12057) );
  INV_X8 U6094 ( .A(n12057), .ZN(n12182) );
  NAND3_X4 U6095 ( .A1(n5287), .A2(n9941), .A3(n5476), .ZN(didKill) );
  INV_X8 U6096 ( .A(net362342), .ZN(net368225) );
  INV_X8 U6097 ( .A(n9680), .ZN(n9722) );
  NOR2_X2 U6098 ( .A1(idOut_114_), .A2(idOut_115_), .ZN(n9979) );
  INV_X4 U6099 ( .A(n10098), .ZN(n5918) );
  INV_X8 U6100 ( .A(n6570), .ZN(n6568) );
  INV_X4 U6101 ( .A(n9766), .ZN(n12944) );
  NOR2_X2 U6102 ( .A1(idOut_25_), .A2(idOut_29_), .ZN(n12945) );
  AOI21_X2 U6103 ( .B1(n6521), .B2(n6523), .A(net368195), .ZN(n11484) );
  NOR2_X2 U6104 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  NOR2_X2 U6105 ( .A1(n7975), .A2(n6531), .ZN(n7980) );
  NOR2_X2 U6106 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  NAND2_X2 U6107 ( .A1(net367029), .A2(net376417), .ZN(n9882) );
  INV_X16 U6108 ( .A(net368787), .ZN(net366911) );
  NOR2_X2 U6109 ( .A1(net366923), .A2(n5550), .ZN(n7704) );
  NOR2_X2 U6110 ( .A1(net366923), .A2(n5531), .ZN(n7699) );
  NOR2_X2 U6111 ( .A1(net366923), .A2(n5533), .ZN(n7720) );
  NOR2_X2 U6112 ( .A1(net366923), .A2(n5536), .ZN(n7729) );
  NOR2_X2 U6113 ( .A1(net366923), .A2(n5548), .ZN(n7689) );
  NOR2_X2 U6114 ( .A1(net366923), .A2(n5546), .ZN(n7683) );
  INV_X1 U6115 ( .A(net361907), .ZN(net377700) );
  NOR2_X2 U6116 ( .A1(net366923), .A2(n5538), .ZN(n7461) );
  NOR2_X2 U6117 ( .A1(net366923), .A2(n5540), .ZN(n7466) );
  NOR2_X2 U6118 ( .A1(net366923), .A2(n5539), .ZN(n7465) );
  NOR2_X2 U6119 ( .A1(n7847), .A2(n7850), .ZN(n7848) );
  AOI21_X2 U6120 ( .B1(n7918), .B2(n7917), .A(net366951), .ZN(n7922) );
  AOI21_X2 U6121 ( .B1(n7914), .B2(n7913), .A(net366925), .ZN(n7915) );
  INV_X4 U6122 ( .A(n11895), .ZN(n11898) );
  NOR2_X1 U6123 ( .A1(n6829), .A2(n8190), .ZN(n8193) );
  NOR2_X1 U6124 ( .A1(n6830), .A2(n6829), .ZN(n8189) );
  NOR2_X1 U6125 ( .A1(n6821), .A2(n8190), .ZN(n8186) );
  NOR2_X2 U6126 ( .A1(n6821), .A2(n6834), .ZN(n8204) );
  NOR2_X2 U6127 ( .A1(n6821), .A2(n6830), .ZN(n8202) );
  NOR2_X1 U6128 ( .A1(n6834), .A2(n6829), .ZN(n8199) );
  OAI21_X1 U6129 ( .B1(n6618), .B2(n6563), .A(n6560), .ZN(n9620) );
  INV_X8 U6130 ( .A(n13533), .ZN(n6532) );
  OAI21_X2 U6131 ( .B1(n8971), .B2(n9049), .A(n9053), .ZN(n8974) );
  INV_X4 U6132 ( .A(n13532), .ZN(n6516) );
  NAND3_X1 U6133 ( .A1(n9196), .A2(n6565), .A3(n5345), .ZN(n9760) );
  OAI21_X2 U6134 ( .B1(n6562), .B2(n9546), .A(n6515), .ZN(n9550) );
  INV_X4 U6135 ( .A(n5714), .ZN(n6556) );
  NAND3_X2 U6136 ( .A1(n13301), .A2(n13335), .A3(n5455), .ZN(n13433) );
  OAI21_X2 U6137 ( .B1(n6562), .B2(n9504), .A(n6523), .ZN(n9508) );
  AOI21_X1 U6138 ( .B1(n9195), .B2(n13527), .A(n9194), .ZN(n9198) );
  NOR2_X1 U6139 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  AOI211_X2 U6140 ( .C1(aluBoi_aluBoi_shft_sraout[1]), .C2(n5460), .A(n13272), 
        .B(net358591), .ZN(n13273) );
  NOR2_X1 U6141 ( .A1(n5387), .A2(n5319), .ZN(net358591) );
  NOR2_X1 U6142 ( .A1(n6569), .A2(n5516), .ZN(n9973) );
  INV_X16 U6143 ( .A(n6506), .ZN(aluBoi_aluBoi_shft_sraout[31]) );
  INV_X8 U6144 ( .A(n13705), .ZN(n6506) );
  OAI21_X1 U6145 ( .B1(n6569), .B2(n5349), .A(idOut_117_), .ZN(n9984) );
  NOR2_X2 U6146 ( .A1(difHold), .A2(n5476), .ZN(n9993) );
  INV_X4 U6147 ( .A(n1205), .ZN(n13673) );
  OAI21_X2 U6148 ( .B1(n13152), .B2(n13151), .A(n13062), .ZN(n13154) );
  OAI21_X2 U6149 ( .B1(n13162), .B2(n13161), .A(n13062), .ZN(n13164) );
  NAND2_X2 U6150 ( .A1(net368215), .A2(net361801), .ZN(n10814) );
  NOR2_X1 U6151 ( .A1(n13706), .A2(net368195), .ZN(n10811) );
  AOI21_X1 U6152 ( .B1(n7761), .B2(n9863), .A(n6531), .ZN(n9864) );
  NOR2_X2 U6153 ( .A1(n11069), .A2(n11068), .ZN(n11074) );
  NOR2_X2 U6154 ( .A1(n10504), .A2(net368209), .ZN(n10505) );
  NOR2_X2 U6155 ( .A1(n6541), .A2(net368209), .ZN(n10698) );
  NOR2_X2 U6156 ( .A1(net368498), .A2(net368209), .ZN(n10484) );
  OAI22_X2 U6157 ( .A1(n11812), .A2(net368467), .B1(n5030), .B2(net368211), 
        .ZN(n11983) );
  NAND3_X2 U6158 ( .A1(n10953), .A2(net361629), .A3(n10952), .ZN(n10937) );
  INV_X2 U6159 ( .A(n6346), .ZN(n7264) );
  INV_X4 U6160 ( .A(n7950), .ZN(n7951) );
  OAI21_X1 U6161 ( .B1(net366921), .B2(n5401), .A(net366967), .ZN(n7445) );
  NAND2_X2 U6162 ( .A1(regBoiz_regfile_31__14_), .A2(net366937), .ZN(n7447) );
  OAI21_X1 U6163 ( .B1(net366921), .B2(n5400), .A(net366967), .ZN(n7435) );
  OAI21_X1 U6164 ( .B1(net366921), .B2(n5399), .A(net366967), .ZN(n7423) );
  OAI21_X1 U6165 ( .B1(net366919), .B2(n5398), .A(net366969), .ZN(n7413) );
  INV_X2 U6166 ( .A(n6295), .ZN(n7024) );
  NOR2_X2 U6167 ( .A1(n7991), .A2(n5444), .ZN(n7992) );
  NAND3_X2 U6168 ( .A1(n5422), .A2(n7980), .A3(n7979), .ZN(n7987) );
  NAND3_X1 U6169 ( .A1(n7984), .A2(n7983), .A3(net366965), .ZN(n7985) );
  NAND3_X2 U6170 ( .A1(net369316), .A2(net366965), .A3(n5959), .ZN(n8005) );
  NOR2_X2 U6171 ( .A1(n8004), .A2(n8003), .ZN(n8011) );
  NOR2_X2 U6172 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  NOR2_X2 U6173 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND3_X2 U6174 ( .A1(net366997), .A2(n5959), .A3(net369316), .ZN(n8018) );
  NAND3_X2 U6175 ( .A1(net366949), .A2(n8015), .A3(net366997), .ZN(n8016) );
  AOI21_X1 U6176 ( .B1(n7784), .B2(n7783), .A(net366951), .ZN(n7788) );
  INV_X4 U6177 ( .A(n6023), .ZN(n7349) );
  AOI22_X1 U6178 ( .A1(regBoiz_regfile_28__12_), .A2(net367003), .B1(
        regBoiz_regfile_30__12_), .B2(net366985), .ZN(n7372) );
  AOI22_X1 U6179 ( .A1(regBoiz_regfile_29__12_), .A2(net367001), .B1(
        regBoiz_regfile_31__12_), .B2(net366985), .ZN(n7371) );
  AOI21_X2 U6180 ( .B1(n7881), .B2(n7880), .A(net366949), .ZN(n7885) );
  AOI21_X2 U6181 ( .B1(n7883), .B2(n7882), .A(net366927), .ZN(n7884) );
  OAI21_X2 U6182 ( .B1(n7871), .B2(n7870), .A(net366999), .ZN(n7879) );
  AOI21_X1 U6183 ( .B1(n7867), .B2(n7866), .A(net366949), .ZN(n7871) );
  AOI21_X1 U6184 ( .B1(n7873), .B2(n7872), .A(net366949), .ZN(n7877) );
  AOI21_X1 U6185 ( .B1(n7875), .B2(n7874), .A(net366927), .ZN(n7876) );
  INV_X4 U6186 ( .A(n11857), .ZN(n6091) );
  NAND2_X2 U6187 ( .A1(n5943), .A2(n12464), .ZN(n12193) );
  NAND3_X2 U6188 ( .A1(n7709), .A2(n7708), .A3(n8147), .ZN(n7718) );
  OAI21_X1 U6189 ( .B1(n5644), .B2(n7704), .A(n6793), .ZN(n7709) );
  NAND3_X2 U6190 ( .A1(n7716), .A2(n7715), .A3(n7714), .ZN(n7717) );
  NOR2_X1 U6191 ( .A1(net369316), .A2(net366997), .ZN(n7714) );
  OAI21_X1 U6192 ( .B1(n7712), .B2(n7711), .A(n6793), .ZN(n7716) );
  NAND3_X2 U6193 ( .A1(n7703), .A2(n7702), .A3(n7701), .ZN(n7719) );
  NOR2_X2 U6194 ( .A1(net366967), .A2(net369316), .ZN(n7701) );
  AOI211_X2 U6195 ( .C1(n7725), .C2(n7724), .A(net364906), .B(net366997), .ZN(
        n7733) );
  AOI211_X2 U6196 ( .C1(n7731), .C2(n7730), .A(net366965), .B(net364906), .ZN(
        n7732) );
  OAI21_X2 U6197 ( .B1(n7728), .B2(n7727), .A(n6793), .ZN(n7731) );
  NAND3_X2 U6198 ( .A1(n7695), .A2(n7694), .A3(n7693), .ZN(n7696) );
  NAND3_X2 U6199 ( .A1(n7688), .A2(n7687), .A3(n7686), .ZN(n7697) );
  NAND3_X1 U6200 ( .A1(n7681), .A2(n7680), .A3(n8144), .ZN(n7698) );
  OAI22_X1 U6201 ( .A1(net375526), .A2(net375527), .B1(net375528), .B2(
        net366989), .ZN(net375525) );
  AOI21_X2 U6202 ( .B1(n7320), .B2(n7319), .A(n7336), .ZN(n7321) );
  NOR2_X1 U6203 ( .A1(net366949), .A2(n7316), .ZN(n7320) );
  NOR3_X2 U6204 ( .A1(n7343), .A2(net366949), .A3(n7342), .ZN(n7344) );
  NOR3_X1 U6205 ( .A1(net366919), .A2(n7343), .A3(n7339), .ZN(n7345) );
  INV_X2 U6206 ( .A(n6457), .ZN(n7071) );
  INV_X2 U6207 ( .A(n6255), .ZN(n7086) );
  NOR2_X2 U6208 ( .A1(net369316), .A2(n8106), .ZN(n8038) );
  AOI22_X2 U6209 ( .A1(n11146), .A2(n5043), .B1(n11144), .B2(n11145), .ZN(
        n11148) );
  INV_X4 U6210 ( .A(n12052), .ZN(n6229) );
  OAI21_X2 U6211 ( .B1(n5641), .B2(n7458), .A(net366967), .ZN(n7459) );
  NOR2_X2 U6212 ( .A1(net366923), .A2(n5526), .ZN(n7458) );
  OAI21_X1 U6213 ( .B1(n5640), .B2(n7457), .A(net367001), .ZN(n7460) );
  NOR2_X2 U6214 ( .A1(net366923), .A2(n5525), .ZN(n7457) );
  OAI21_X2 U6215 ( .B1(n5431), .B2(n7491), .A(net366967), .ZN(n7492) );
  OAI21_X2 U6216 ( .B1(n5437), .B2(n7487), .A(net366967), .ZN(n7488) );
  OAI21_X1 U6217 ( .B1(n5427), .B2(n7469), .A(net367001), .ZN(n7472) );
  OAI21_X2 U6218 ( .B1(n5432), .B2(n7461), .A(net367001), .ZN(n7464) );
  OAI21_X1 U6219 ( .B1(n5642), .B2(n7462), .A(net366967), .ZN(n7463) );
  OAI21_X2 U6220 ( .B1(n5643), .B2(n7465), .A(net367001), .ZN(n7468) );
  OAI21_X2 U6221 ( .B1(n5433), .B2(n7466), .A(net366967), .ZN(n7467) );
  AOI21_X2 U6222 ( .B1(n7615), .B2(n7614), .A(net366999), .ZN(n7623) );
  AOI21_X2 U6223 ( .B1(n7826), .B2(n7825), .A(net366925), .ZN(n7827) );
  NAND3_X1 U6224 ( .A1(n7816), .A2(net366997), .A3(n5959), .ZN(n7832) );
  NAND3_X1 U6225 ( .A1(n7814), .A2(net365293), .A3(net366965), .ZN(n7833) );
  NAND3_X1 U6226 ( .A1(n7839), .A2(net366947), .A3(n5333), .ZN(n7844) );
  NAND3_X1 U6227 ( .A1(n7842), .A2(net366947), .A3(n7841), .ZN(n7843) );
  NAND3_X1 U6228 ( .A1(n7837), .A2(n5333), .A3(net366919), .ZN(n7845) );
  NAND3_X1 U6229 ( .A1(n7835), .A2(n7841), .A3(net366919), .ZN(n7846) );
  NAND3_X1 U6230 ( .A1(n7810), .A2(n5959), .A3(net366965), .ZN(n7811) );
  NAND3_X1 U6231 ( .A1(n7808), .A2(net366997), .A3(net365293), .ZN(n7812) );
  NAND3_X1 U6232 ( .A1(net366919), .A2(n7852), .A3(n7851), .ZN(n7859) );
  NAND3_X1 U6233 ( .A1(n7855), .A2(n7854), .A3(net366919), .ZN(n7858) );
  AOI21_X2 U6234 ( .B1(n7904), .B2(n7903), .A(net366951), .ZN(n7908) );
  AOI21_X2 U6235 ( .B1(n7906), .B2(n7905), .A(net366925), .ZN(n7907) );
  AOI21_X2 U6236 ( .B1(n7898), .B2(n7897), .A(net366951), .ZN(n7902) );
  AOI21_X2 U6237 ( .B1(n7900), .B2(n7899), .A(net366925), .ZN(n7901) );
  AOI21_X2 U6238 ( .B1(n7912), .B2(n7911), .A(net366951), .ZN(n7916) );
  NAND3_X2 U6239 ( .A1(n12364), .A2(n12562), .A3(n12363), .ZN(n12365) );
  INV_X4 U6240 ( .A(net359876), .ZN(net368461) );
  NAND2_X2 U6241 ( .A1(aluBoi_multOut[0]), .A2(n5319), .ZN(net359876) );
  NAND2_X2 U6242 ( .A1(net376602), .A2(n6055), .ZN(n8880) );
  OAI21_X2 U6243 ( .B1(n9474), .B2(n9473), .A(n8884), .ZN(n9462) );
  OAI21_X2 U6244 ( .B1(n9464), .B2(n9465), .A(n9463), .ZN(n8764) );
  INV_X4 U6245 ( .A(n9076), .ZN(n8623) );
  NOR2_X2 U6246 ( .A1(n6613), .A2(n9682), .ZN(n9683) );
  NAND2_X2 U6247 ( .A1(daddr[13]), .A2(net368221), .ZN(n9834) );
  AOI21_X2 U6248 ( .B1(n8079), .B2(n8078), .A(net366967), .ZN(n8082) );
  AOI21_X2 U6249 ( .B1(n8076), .B2(n8075), .A(net366999), .ZN(n8084) );
  AOI21_X1 U6250 ( .B1(n8096), .B2(n8095), .A(net366951), .ZN(n8100) );
  OAI21_X2 U6251 ( .B1(n8094), .B2(n8093), .A(net366999), .ZN(n8102) );
  AOI21_X1 U6252 ( .B1(n8090), .B2(n8089), .A(net366951), .ZN(n8094) );
  NOR3_X2 U6253 ( .A1(net366965), .A2(n8104), .A3(n8106), .ZN(net364898) );
  AOI21_X2 U6254 ( .B1(n8108), .B2(n8107), .A(net366951), .ZN(n8112) );
  AOI21_X2 U6255 ( .B1(n8114), .B2(n8113), .A(net366951), .ZN(n8118) );
  AOI21_X2 U6256 ( .B1(n8116), .B2(n8115), .A(net366925), .ZN(n8117) );
  NOR3_X2 U6257 ( .A1(n8153), .A2(n5587), .A3(n8152), .ZN(n8154) );
  NOR3_X2 U6258 ( .A1(n8151), .A2(n5586), .A3(n8150), .ZN(n8155) );
  NAND3_X2 U6259 ( .A1(n8147), .A2(n8146), .A3(n8145), .ZN(n8148) );
  AOI21_X2 U6260 ( .B1(n9665), .B2(n6560), .A(n9664), .ZN(n9668) );
  OAI21_X2 U6261 ( .B1(n9641), .B2(n10850), .A(n9640), .ZN(n12983) );
  NOR2_X2 U6262 ( .A1(n6562), .A2(n9638), .ZN(n9641) );
  OAI21_X2 U6263 ( .B1(n9619), .B2(net361631), .A(n9618), .ZN(n12960) );
  NOR2_X2 U6264 ( .A1(n6562), .A2(n9616), .ZN(n9619) );
  OAI21_X2 U6265 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n13085) );
  NOR2_X2 U6266 ( .A1(n6562), .A2(n9652), .ZN(n9656) );
  AOI21_X1 U6267 ( .B1(n9672), .B2(n6560), .A(n9671), .ZN(n9675) );
  NAND3_X2 U6268 ( .A1(n12151), .A2(n12150), .A3(aluBoi_multBoi_temppp[57]), 
        .ZN(net359767) );
  NOR2_X1 U6269 ( .A1(n6569), .A2(n5513), .ZN(n9966) );
  NOR2_X1 U6270 ( .A1(n6569), .A2(n5517), .ZN(n9976) );
  OAI21_X2 U6271 ( .B1(n5347), .B2(n10332), .A(n6548), .ZN(n10344) );
  NAND3_X2 U6272 ( .A1(n13321), .A2(n5455), .A3(n13493), .ZN(n9994) );
  NOR3_X2 U6273 ( .A1(n8708), .A2(n8223), .A3(n8222), .ZN(n8224) );
  NAND3_X2 U6274 ( .A1(n8196), .A2(n8195), .A3(n8194), .ZN(n8226) );
  NOR2_X2 U6275 ( .A1(n5353), .A2(n5318), .ZN(n1209) );
  NOR2_X2 U6276 ( .A1(n5511), .A2(wbRwh[1]), .ZN(n99) );
  NOR2_X2 U6277 ( .A1(wbRwh[0]), .A2(wbRwh[1]), .ZN(n134) );
  OAI21_X2 U6278 ( .B1(n9496), .B2(n10346), .A(n9495), .ZN(n12975) );
  NOR2_X2 U6279 ( .A1(n6562), .A2(n9493), .ZN(n9496) );
  OAI21_X2 U6280 ( .B1(n6562), .B2(n9621), .A(n6618), .ZN(n9622) );
  OAI21_X2 U6281 ( .B1(n9614), .B2(n10575), .A(n9613), .ZN(n13042) );
  NOR2_X2 U6282 ( .A1(n6562), .A2(n9611), .ZN(n9614) );
  INV_X4 U6283 ( .A(n13535), .ZN(n6524) );
  OAI21_X1 U6284 ( .B1(n6525), .B2(n6564), .A(n6561), .ZN(n9517) );
  OAI21_X1 U6285 ( .B1(n6527), .B2(n6563), .A(n6560), .ZN(n9602) );
  OAI21_X2 U6286 ( .B1(n6562), .B2(n9498), .A(n6521), .ZN(n9502) );
  OAI21_X2 U6287 ( .B1(n6562), .B2(n9552), .A(net368572), .ZN(n9556) );
  OAI21_X2 U6288 ( .B1(n6562), .B2(n9537), .A(n6517), .ZN(n9541) );
  OAI21_X1 U6289 ( .B1(n6562), .B2(n9559), .A(n5309), .ZN(n9563) );
  NAND3_X2 U6290 ( .A1(n9599), .A2(n9598), .A3(n9597), .ZN(n13237) );
  INV_X4 U6291 ( .A(n9760), .ZN(n12940) );
  INV_X2 U6292 ( .A(n5758), .ZN(n8316) );
  NAND3_X2 U6293 ( .A1(n13342), .A2(n13499), .A3(n13341), .ZN(n13356) );
  NOR2_X2 U6294 ( .A1(n5312), .A2(n5343), .ZN(n13341) );
  NOR2_X2 U6295 ( .A1(n5312), .A2(n13340), .ZN(n13307) );
  INV_X16 U6296 ( .A(n6580), .ZN(n6585) );
  OAI21_X2 U6297 ( .B1(n6562), .B2(n9589), .A(n6529), .ZN(n9593) );
  NOR2_X2 U6298 ( .A1(n6611), .A2(n5484), .ZN(n12943) );
  NOR2_X1 U6299 ( .A1(n12666), .A2(n6551), .ZN(n10078) );
  NOR2_X2 U6300 ( .A1(n6569), .A2(n5515), .ZN(n9971) );
  NOR2_X2 U6301 ( .A1(n12053), .A2(n6573), .ZN(n10067) );
  NOR2_X2 U6302 ( .A1(n12054), .A2(n6573), .ZN(n10053) );
  NOR2_X1 U6303 ( .A1(n12681), .A2(n6551), .ZN(n10092) );
  NOR2_X2 U6304 ( .A1(n10089), .A2(n6573), .ZN(n10094) );
  NOR2_X2 U6305 ( .A1(n12833), .A2(n10345), .ZN(n10300) );
  NOR2_X1 U6306 ( .A1(n10850), .A2(n6574), .ZN(n10293) );
  NOR2_X1 U6307 ( .A1(net362485), .A2(n6574), .ZN(n10361) );
  INV_X8 U6308 ( .A(n13710), .ZN(n6617) );
  NAND3_X1 U6309 ( .A1(n8261), .A2(n8697), .A3(n8698), .ZN(n13710) );
  NAND3_X2 U6310 ( .A1(n8801), .A2(n8800), .A3(n8799), .ZN(n10422) );
  NAND3_X2 U6311 ( .A1(n8921), .A2(n5457), .A3(n8920), .ZN(n10424) );
  NAND3_X2 U6312 ( .A1(n8868), .A2(n5457), .A3(n8867), .ZN(n10425) );
  NAND3_X1 U6313 ( .A1(n9721), .A2(n5457), .A3(n9720), .ZN(n10497) );
  NOR2_X1 U6314 ( .A1(n11669), .A2(n5335), .ZN(n11437) );
  INV_X4 U6315 ( .A(n1146), .ZN(n13712) );
  NOR2_X1 U6316 ( .A1(n12876), .A2(n5509), .ZN(n12875) );
  NAND3_X2 U6317 ( .A1(ifInst[31]), .A2(n13491), .A3(n5455), .ZN(n12917) );
  NAND3_X2 U6318 ( .A1(ifInst[31]), .A2(n5455), .A3(n13493), .ZN(n13324) );
  NAND3_X1 U6319 ( .A1(ifInst[28]), .A2(n13491), .A3(n12921), .ZN(n13322) );
  NOR2_X2 U6320 ( .A1(ifInst[30]), .A2(ifInst[29]), .ZN(n12921) );
  AOI222_X2 U6321 ( .A1(n13019), .A2(n13141), .B1(aluBoi_multBoi_temppp[18]), 
        .B2(net368069), .C1(n5316), .C2(aluBoi_imm32w_5_), .ZN(n13146) );
  NOR2_X2 U6322 ( .A1(idOut_25_), .A2(didMult), .ZN(n12939) );
  OAI21_X2 U6323 ( .B1(n13238), .B2(n13237), .A(n6605), .ZN(n13241) );
  NOR2_X1 U6324 ( .A1(n5387), .A2(n5471), .ZN(net358618) );
  AOI211_X2 U6325 ( .C1(aluBoi_aluBoi_shft_sraout[2]), .C2(n5460), .A(n13261), 
        .B(net358604), .ZN(n13262) );
  NOR2_X1 U6326 ( .A1(n5387), .A2(n5304), .ZN(net358604) );
  NAND3_X2 U6327 ( .A1(n5575), .A2(n13293), .A3(n13292), .ZN(n13294) );
  NAND3_X2 U6328 ( .A1(n13289), .A2(ifInst[1]), .A3(n5459), .ZN(n13293) );
  AOI21_X2 U6329 ( .B1(n13291), .B2(n5343), .A(n5555), .ZN(n13292) );
  NOR2_X2 U6330 ( .A1(ifInst[31]), .A2(ifInst[29]), .ZN(n13301) );
  NOR3_X2 U6331 ( .A1(n13326), .A2(n6586), .A3(n5474), .ZN(n13327) );
  NOR2_X1 U6332 ( .A1(ifInst[1]), .A2(ifInst[3]), .ZN(n13319) );
  NOR2_X2 U6333 ( .A1(n5312), .A2(n5456), .ZN(n13317) );
  NOR2_X2 U6334 ( .A1(n5343), .A2(n13340), .ZN(n13334) );
  NAND3_X2 U6335 ( .A1(ifInst[29]), .A2(ifInst[30]), .A3(n13497), .ZN(n13358)
         );
  OAI21_X2 U6336 ( .B1(n13499), .B2(n13357), .A(n13356), .ZN(n13348) );
  NAND3_X2 U6337 ( .A1(ifInst[29]), .A2(n5455), .A3(n13497), .ZN(n13400) );
  OAI21_X2 U6338 ( .B1(n5689), .B2(n6611), .A(n3354), .ZN(n4799) );
  NAND3_X2 U6339 ( .A1(n9947), .A2(n9946), .A3(n9945), .ZN(n9999) );
  OAI21_X2 U6340 ( .B1(n10004), .B2(n10003), .A(n10408), .ZN(n10017) );
  INV_X4 U6341 ( .A(n6944), .ZN(n6943) );
  NOR3_X1 U6342 ( .A1(net368502), .A2(n10916), .A3(n10915), .ZN(n10920) );
  NAND2_X2 U6343 ( .A1(n10890), .A2(n11232), .ZN(n10895) );
  OAI21_X2 U6344 ( .B1(n9869), .B2(net363057), .A(n9875), .ZN(n9870) );
  NAND2_X2 U6345 ( .A1(n10949), .A2(net368201), .ZN(n6439) );
  NOR2_X1 U6346 ( .A1(net368519), .A2(net368195), .ZN(n10810) );
  NOR2_X2 U6347 ( .A1(n6432), .A2(n11049), .ZN(n11013) );
  NOR3_X2 U6348 ( .A1(n9837), .A2(n9836), .A3(n9835), .ZN(n9838) );
  NOR2_X2 U6349 ( .A1(net368498), .A2(net368203), .ZN(net362255) );
  INV_X4 U6350 ( .A(net359986), .ZN(net368445) );
  OAI21_X1 U6351 ( .B1(n10941), .B2(n10945), .A(n10964), .ZN(n10946) );
  NAND2_X2 U6352 ( .A1(n5774), .A2(n5775), .ZN(net375304) );
  NOR2_X2 U6353 ( .A1(net368195), .A2(n13706), .ZN(n10775) );
  NAND3_X2 U6354 ( .A1(net366997), .A2(n7935), .A3(net366919), .ZN(n7936) );
  INV_X4 U6355 ( .A(n11576), .ZN(n11658) );
  AOI21_X2 U6356 ( .B1(n11614), .B2(n5893), .A(n11543), .ZN(n11569) );
  INV_X4 U6357 ( .A(n11412), .ZN(n11415) );
  OAI21_X2 U6358 ( .B1(n11828), .B2(n11827), .A(n11799), .ZN(n11803) );
  INV_X4 U6359 ( .A(n10578), .ZN(n10552) );
  INV_X4 U6360 ( .A(n6039), .ZN(n6040) );
  NOR2_X2 U6361 ( .A1(n10956), .A2(n10843), .ZN(n10715) );
  NAND2_X2 U6362 ( .A1(aluBoi_multOut[1]), .A2(n5304), .ZN(net359986) );
  OAI22_X2 U6363 ( .A1(net361801), .A2(net368439), .B1(net368185), .B2(
        net362124), .ZN(net362140) );
  NAND2_X2 U6364 ( .A1(n11504), .A2(n11577), .ZN(n11505) );
  NOR2_X2 U6365 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  INV_X16 U6366 ( .A(net368191), .ZN(net368187) );
  NAND2_X2 U6367 ( .A1(n6165), .A2(n6166), .ZN(n9881) );
  NOR2_X2 U6368 ( .A1(n8628), .A2(n9104), .ZN(n8722) );
  OAI21_X2 U6369 ( .B1(n11874), .B2(n11873), .A(n11872), .ZN(n11880) );
  INV_X4 U6370 ( .A(n12435), .ZN(n12078) );
  OAI21_X2 U6371 ( .B1(n5990), .B2(n11260), .A(n11259), .ZN(n11335) );
  INV_X4 U6372 ( .A(net360631), .ZN(n5787) );
  AOI21_X2 U6373 ( .B1(n12178), .B2(n12256), .A(n12177), .ZN(n12179) );
  INV_X4 U6374 ( .A(n12260), .ZN(n12265) );
  NOR2_X2 U6375 ( .A1(n7745), .A2(n9848), .ZN(n7753) );
  NOR3_X1 U6376 ( .A1(n7758), .A2(net366919), .A3(net369316), .ZN(n7763) );
  INV_X16 U6377 ( .A(net369143), .ZN(net369158) );
  INV_X4 U6378 ( .A(net361832), .ZN(net376826) );
  INV_X8 U6379 ( .A(n6426), .ZN(n6427) );
  INV_X4 U6380 ( .A(n11156), .ZN(n6426) );
  INV_X4 U6381 ( .A(n11051), .ZN(n6530) );
  NOR2_X1 U6382 ( .A1(aluBoi_aluBoi_shft_sllout[10]), .A2(
        aluBoi_aluBoi_shft_sllout[11]), .ZN(n8363) );
  NOR2_X1 U6383 ( .A1(aluBoi_aluBoi_shft_sraout[11]), .A2(
        aluBoi_aluBoi_shft_sraout[10]), .ZN(n8377) );
  NOR2_X1 U6384 ( .A1(aluBoi_aluBoi_shft_sraout[17]), .A2(
        aluBoi_aluBoi_shft_sraout[16]), .ZN(n8375) );
  NOR3_X1 U6385 ( .A1(aluBoi_aluBoi_shft_sraout[6]), .A2(
        aluBoi_aluBoi_shft_sraout[8]), .A3(aluBoi_aluBoi_shft_sraout[7]), .ZN(
        n8369) );
  NOR2_X1 U6386 ( .A1(aluBoi_aluBoi_shft_sraout[4]), .A2(
        aluBoi_aluBoi_shft_sraout[3]), .ZN(n8367) );
  NOR3_X1 U6387 ( .A1(aluBoi_aluBoi_shft_sllout[0]), .A2(
        aluBoi_aluBoi_shft_sllout[2]), .A3(aluBoi_aluBoi_shft_sllout[1]), .ZN(
        n8357) );
  INV_X16 U6388 ( .A(n5388), .ZN(net368217) );
  INV_X4 U6389 ( .A(net359601), .ZN(net368183) );
  NAND3_X1 U6390 ( .A1(n12054), .A2(n12053), .A3(n12060), .ZN(n12056) );
  INV_X4 U6391 ( .A(net359754), .ZN(net368435) );
  NAND2_X2 U6392 ( .A1(aluBoi_multOut[2]), .A2(n5471), .ZN(net359754) );
  INV_X8 U6393 ( .A(net368439), .ZN(net359752) );
  AOI21_X1 U6394 ( .B1(n12460), .B2(n12573), .A(n12570), .ZN(n12462) );
  NOR3_X1 U6395 ( .A1(n9866), .A2(net369316), .A3(n9848), .ZN(n7742) );
  NOR2_X2 U6396 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  NAND3_X2 U6397 ( .A1(n7323), .A2(n7322), .A3(n7321), .ZN(n7348) );
  INV_X16 U6398 ( .A(net369148), .ZN(net369248) );
  BUF_X4 U6399 ( .A(net369138), .Z(net369139) );
  NAND3_X2 U6400 ( .A1(n9461), .A2(n8935), .A3(n8934), .ZN(n9052) );
  OAI21_X1 U6401 ( .B1(n13706), .B2(n6563), .A(n6560), .ZN(n9639) );
  OAI21_X1 U6402 ( .B1(net368519), .B2(n6563), .A(n6560), .ZN(n9617) );
  OAI21_X1 U6403 ( .B1(n6539), .B2(n6563), .A(n6560), .ZN(n9653) );
  NOR2_X2 U6404 ( .A1(n11692), .A2(n11955), .ZN(n11693) );
  NOR2_X2 U6405 ( .A1(n10805), .A2(n5043), .ZN(n10808) );
  INV_X1 U6406 ( .A(n6568), .ZN(n5756) );
  INV_X4 U6407 ( .A(n10190), .ZN(n5757) );
  NAND3_X2 U6408 ( .A1(n7460), .A2(n7459), .A3(net365399), .ZN(n7476) );
  NAND3_X2 U6409 ( .A1(n9544), .A2(n9543), .A3(n9542), .ZN(n9557) );
  NOR3_X1 U6410 ( .A1(n13124), .A2(n13237), .A3(n13113), .ZN(n9606) );
  NOR3_X2 U6411 ( .A1(n8378), .A2(n5717), .A3(n5393), .ZN(n8379) );
  NAND3_X2 U6412 ( .A1(n8377), .A2(n8376), .A3(n8375), .ZN(n8378) );
  NOR2_X2 U6413 ( .A1(n8374), .A2(n8373), .ZN(n8380) );
  NAND3_X2 U6414 ( .A1(n8369), .A2(n8368), .A3(n8367), .ZN(n8374) );
  NAND3_X2 U6415 ( .A1(n8372), .A2(n8371), .A3(n8370), .ZN(n8373) );
  NOR3_X1 U6416 ( .A1(n8359), .A2(aluBoi_aluBoi_shft_sllout[6]), .A3(
        aluBoi_aluBoi_shft_sllout[5]), .ZN(n8366) );
  NAND3_X2 U6417 ( .A1(n8358), .A2(n8357), .A3(n8356), .ZN(n8359) );
  NOR2_X1 U6418 ( .A1(aluBoi_aluBoi_shft_sllout[4]), .A2(
        aluBoi_aluBoi_shft_sllout[3]), .ZN(n8358) );
  NOR2_X1 U6419 ( .A1(aluBoi_aluBoi_shft_sllout[8]), .A2(
        aluBoi_aluBoi_shft_sllout[7]), .ZN(n8356) );
  NOR3_X2 U6420 ( .A1(n9111), .A2(n9110), .A3(n9109), .ZN(n9112) );
  NAND3_X1 U6421 ( .A1(n13083), .A2(n12958), .A3(n12980), .ZN(n9111) );
  NOR3_X2 U6422 ( .A1(n9048), .A2(n9047), .A3(n9046), .ZN(n9114) );
  NOR2_X1 U6423 ( .A1(n13091), .A2(n9063), .ZN(n9113) );
  OAI21_X2 U6424 ( .B1(n9476), .B2(n9475), .A(n13220), .ZN(n9481) );
  NAND3_X1 U6425 ( .A1(n13071), .A2(n13059), .A3(n13047), .ZN(n9475) );
  AOI21_X2 U6426 ( .B1(n9478), .B2(n9477), .A(n9766), .ZN(n9479) );
  NOR2_X1 U6427 ( .A1(aluBoi_aluBoi_shft_sraout[15]), .A2(
        aluBoi_aluBoi_shft_sraout[14]), .ZN(n9477) );
  NOR2_X1 U6428 ( .A1(aluBoi_aluBoi_shft_sraout[13]), .A2(
        aluBoi_aluBoi_shft_sraout[12]), .ZN(n9478) );
  AOI21_X2 U6429 ( .B1(n9459), .B2(n9458), .A(n9760), .ZN(n9460) );
  NOR2_X1 U6430 ( .A1(aluBoi_aluBoi_shft_sllout[15]), .A2(
        aluBoi_aluBoi_shft_sllout[14]), .ZN(n9458) );
  NOR2_X1 U6431 ( .A1(aluBoi_aluBoi_shft_sllout[13]), .A2(
        aluBoi_aluBoi_shft_sllout[12]), .ZN(n9459) );
  INV_X2 U6432 ( .A(n11662), .ZN(n6086) );
  INV_X4 U6433 ( .A(net359966), .ZN(net368466) );
  INV_X16 U6434 ( .A(net368183), .ZN(net368179) );
  NAND3_X2 U6435 ( .A1(n12563), .A2(n12565), .A3(n12562), .ZN(n12476) );
  NOR2_X2 U6436 ( .A1(wbRwh[2]), .A2(wbRwh[3]), .ZN(n907) );
  NOR2_X2 U6437 ( .A1(n5565), .A2(wbRwh[4]), .ZN(n271) );
  NOR2_X2 U6438 ( .A1(n5482), .A2(wbRwh[3]), .ZN(n270) );
  OAI21_X1 U6439 ( .B1(n6545), .B2(n6564), .A(n6561), .ZN(n9494) );
  OAI21_X1 U6440 ( .B1(n6541), .B2(n6563), .A(n6560), .ZN(n9633) );
  OAI21_X1 U6441 ( .B1(n6543), .B2(n6563), .A(n6560), .ZN(n9612) );
  OAI21_X1 U6442 ( .B1(n6521), .B2(n6564), .A(n6561), .ZN(n9499) );
  INV_X1 U6443 ( .A(n9200), .ZN(n5728) );
  OAI21_X1 U6444 ( .B1(n5309), .B2(n6564), .A(n6561), .ZN(n9560) );
  OAI21_X2 U6445 ( .B1(n6509), .B2(n6564), .A(n6561), .ZN(n9578) );
  INV_X8 U6446 ( .A(n6815), .ZN(n6808) );
  NOR3_X1 U6447 ( .A1(ifInst[25]), .A2(ifInst[6]), .A3(ifInst[4]), .ZN(n2011)
         );
  NOR2_X1 U6448 ( .A1(ifInst[9]), .A2(ifInst[10]), .ZN(n13313) );
  NOR2_X1 U6449 ( .A1(ifInst[7]), .A2(ifInst[8]), .ZN(n13314) );
  OAI21_X1 U6450 ( .B1(n6529), .B2(n6563), .A(n6561), .ZN(n9590) );
  OAI21_X1 U6451 ( .B1(n6523), .B2(n6564), .A(n6561), .ZN(n9505) );
  AOI21_X1 U6452 ( .B1(n5288), .B2(n11316), .A(n6562), .ZN(n9192) );
  AOI21_X1 U6453 ( .B1(n9466), .B2(n9465), .A(n9464), .ZN(n9467) );
  INV_X4 U6454 ( .A(net378052), .ZN(n5856) );
  NAND2_X2 U6455 ( .A1(aluBoi_multBoi_temppp[39]), .A2(net378052), .ZN(
        net361296) );
  OAI21_X2 U6456 ( .B1(n10045), .B2(n9978), .A(n6569), .ZN(n9980) );
  NAND3_X2 U6457 ( .A1(n5916), .A2(n9982), .A3(n5349), .ZN(n10008) );
  INV_X4 U6458 ( .A(n10164), .ZN(n5751) );
  INV_X16 U6459 ( .A(n6534), .ZN(n6535) );
  INV_X8 U6460 ( .A(n13531), .ZN(n6534) );
  OAI21_X1 U6461 ( .B1(n8100), .B2(n8099), .A(net366969), .ZN(n8101) );
  NOR3_X2 U6462 ( .A1(n8126), .A2(n8125), .A3(n8124), .ZN(net364875) );
  NOR3_X1 U6463 ( .A1(n13513), .A2(n9733), .A3(n9732), .ZN(n9781) );
  NAND3_X2 U6464 ( .A1(n13509), .A2(n13510), .A3(n13511), .ZN(n9732) );
  NOR2_X2 U6465 ( .A1(n9557), .A2(n5718), .ZN(n9609) );
  NOR2_X1 U6466 ( .A1(n13181), .A2(n13161), .ZN(n9608) );
  NOR3_X1 U6467 ( .A1(n13259), .A2(n13224), .A3(n13270), .ZN(n9607) );
  NOR3_X1 U6468 ( .A1(n13020), .A2(n13031), .A3(n12983), .ZN(n9642) );
  NOR3_X1 U6469 ( .A1(n13042), .A2(n12960), .A3(n13012), .ZN(n9643) );
  NAND3_X2 U6470 ( .A1(n9523), .A2(n9522), .A3(n9521), .ZN(n9646) );
  NOR2_X1 U6471 ( .A1(n13250), .A2(n13102), .ZN(n9521) );
  NOR3_X1 U6472 ( .A1(n13142), .A2(n12975), .A3(n13131), .ZN(n9523) );
  NOR3_X1 U6473 ( .A1(n13050), .A2(n13283), .A3(n9734), .ZN(n9774) );
  NOR3_X1 U6474 ( .A1(n13085), .A2(n13061), .A3(n13074), .ZN(n9775) );
  AOI21_X2 U6475 ( .B1(n12940), .B2(n8382), .A(n8381), .ZN(n9650) );
  AOI21_X2 U6476 ( .B1(n8380), .B2(n8379), .A(n9766), .ZN(n8381) );
  NOR3_X2 U6477 ( .A1(n5719), .A2(n8364), .A3(n5394), .ZN(n8365) );
  AOI21_X2 U6478 ( .B1(n13220), .B2(n9208), .A(n9207), .ZN(n9649) );
  NAND3_X2 U6479 ( .A1(n9206), .A2(n9205), .A3(n9204), .ZN(n9207) );
  NAND3_X2 U6480 ( .A1(n9114), .A2(n9113), .A3(n9112), .ZN(n9208) );
  NOR3_X2 U6481 ( .A1(n9485), .A2(n9484), .A3(n9483), .ZN(n9648) );
  NAND3_X2 U6482 ( .A1(n9482), .A2(n9481), .A3(n9480), .ZN(n9483) );
  NOR2_X2 U6483 ( .A1(n13222), .A2(n9457), .ZN(n9484) );
  INV_X8 U6484 ( .A(n13708), .ZN(n6613) );
  NAND3_X1 U6485 ( .A1(n8355), .A2(n8709), .A3(n8710), .ZN(n13708) );
  NAND2_X2 U6486 ( .A1(aluBoi_imm32w_3_), .A2(n6556), .ZN(n8697) );
  INV_X4 U6487 ( .A(n9719), .ZN(n6546) );
  INV_X4 U6488 ( .A(n8227), .ZN(n9719) );
  NOR2_X2 U6489 ( .A1(n12540), .A2(net359465), .ZN(n12542) );
  NOR2_X2 U6490 ( .A1(n12581), .A2(n12580), .ZN(n12572) );
  NOR2_X2 U6491 ( .A1(n12575), .A2(n12574), .ZN(n12576) );
  NOR2_X2 U6492 ( .A1(n5318), .A2(dSize[1]), .ZN(n1208) );
  INV_X16 U6493 ( .A(n6828), .ZN(n6826) );
  OAI211_X2 U6494 ( .C1(n9187), .C2(n13222), .A(n9186), .B(n9185), .ZN(n13162)
         );
  OAI21_X2 U6495 ( .B1(n6513), .B2(n6564), .A(n6561), .ZN(n9532) );
  NOR2_X2 U6496 ( .A1(n13290), .A2(n13340), .ZN(n13291) );
  NOR2_X1 U6497 ( .A1(ifInst[3]), .A2(ifInst[4]), .ZN(n13288) );
  NAND3_X1 U6498 ( .A1(n13333), .A2(ifInst[5]), .A3(n5456), .ZN(n13340) );
  NOR2_X1 U6499 ( .A1(ifInst[27]), .A2(ifInst[26]), .ZN(n13335) );
  NAND3_X1 U6500 ( .A1(n8220), .A2(n6816), .A3(n8215), .ZN(n12926) );
  NOR2_X2 U6501 ( .A1(net369164), .A2(n6821), .ZN(n8215) );
  INV_X4 U6502 ( .A(n9779), .ZN(n5768) );
  NOR2_X2 U6503 ( .A1(n10101), .A2(n6573), .ZN(n10106) );
  NOR2_X1 U6504 ( .A1(n10140), .A2(n10139), .ZN(n10141) );
  NOR2_X1 U6505 ( .A1(n10136), .A2(n6577), .ZN(n10142) );
  NAND3_X2 U6506 ( .A1(ifOut_93_), .A2(ifOut_92_), .A3(n10019), .ZN(n10028) );
  AOI21_X2 U6507 ( .B1(n10022), .B2(n10023), .A(n10139), .ZN(n10026) );
  NOR2_X2 U6508 ( .A1(ifOut_92_), .A2(ifOut_93_), .ZN(n10022) );
  NAND3_X2 U6509 ( .A1(ifOut_93_), .A2(n5466), .A3(n10024), .ZN(n10025) );
  NAND3_X1 U6510 ( .A1(ifOut_92_), .A2(n5458), .A3(n10020), .ZN(n10027) );
  NOR2_X2 U6511 ( .A1(n12249), .A2(n6573), .ZN(n10039) );
  NOR2_X2 U6512 ( .A1(n5048), .A2(net359904), .ZN(n12228) );
  NOR2_X1 U6513 ( .A1(n5387), .A2(n5307), .ZN(net358577) );
  NOR3_X1 U6514 ( .A1(idOut_25_), .A2(n5314), .A3(n13281), .ZN(n13282) );
  NOR2_X1 U6515 ( .A1(ifInst[28]), .A2(n13433), .ZN(n13333) );
  NOR2_X2 U6516 ( .A1(n6569), .A2(n5514), .ZN(n9969) );
  NOR2_X1 U6517 ( .A1(n11487), .A2(n6573), .ZN(n10153) );
  NOR2_X2 U6518 ( .A1(n10177), .A2(n6573), .ZN(n10178) );
  NOR2_X1 U6519 ( .A1(n11067), .A2(n6574), .ZN(n10231) );
  NOR2_X1 U6520 ( .A1(n6536), .A2(n6574), .ZN(n10256) );
  AOI21_X1 U6521 ( .B1(n10286), .B2(n10285), .A(n10344), .ZN(n10287) );
  NOR2_X1 U6522 ( .A1(net361808), .A2(n6574), .ZN(n10281) );
  NOR2_X1 U6523 ( .A1(n10309), .A2(n6574), .ZN(n10310) );
  NOR2_X2 U6524 ( .A1(n10333), .A2(n10344), .ZN(n10334) );
  NOR2_X2 U6525 ( .A1(n9777), .A2(n9776), .ZN(n13538) );
  NOR3_X2 U6526 ( .A1(n9646), .A2(n9645), .A3(n9644), .ZN(n9647) );
  OAI21_X2 U6527 ( .B1(n13538), .B2(n5391), .A(n5715), .ZN(n2847) );
  INV_X8 U6528 ( .A(n5317), .ZN(n6606) );
  NAND3_X2 U6529 ( .A1(n8621), .A2(n8620), .A3(n8619), .ZN(n10413) );
  INV_X8 U6530 ( .A(n13711), .ZN(n6619) );
  NAND3_X2 U6531 ( .A1(n8230), .A2(n8229), .A3(n8228), .ZN(n13711) );
  NAND3_X2 U6532 ( .A1(n8551), .A2(n8550), .A3(n8549), .ZN(n10414) );
  NAND3_X2 U6533 ( .A1(n8483), .A2(n8482), .A3(n8481), .ZN(n10417) );
  NAND3_X2 U6534 ( .A1(n8415), .A2(n8414), .A3(n8413), .ZN(n10418) );
  NAND3_X2 U6535 ( .A1(n8448), .A2(n8447), .A3(n8446), .ZN(n10419) );
  NAND3_X2 U6536 ( .A1(n8760), .A2(n8759), .A3(n8758), .ZN(n10420) );
  NAND3_X2 U6537 ( .A1(n8517), .A2(n8516), .A3(n8515), .ZN(n10421) );
  NAND3_X2 U6538 ( .A1(n8969), .A2(n5457), .A3(n8968), .ZN(n10423) );
  NAND3_X2 U6539 ( .A1(n8836), .A2(n5457), .A3(n8835), .ZN(n10426) );
  NAND3_X2 U6540 ( .A1(n9007), .A2(n5457), .A3(n9006), .ZN(n10427) );
  NAND3_X2 U6541 ( .A1(n9041), .A2(n5457), .A3(n9040), .ZN(n10428) );
  NAND3_X2 U6542 ( .A1(n9149), .A2(n5457), .A3(n9148), .ZN(n10429) );
  NAND3_X1 U6543 ( .A1(n9183), .A2(n5457), .A3(n9182), .ZN(n10430) );
  NAND3_X1 U6544 ( .A1(n9340), .A2(n5457), .A3(n9339), .ZN(n10431) );
  NAND3_X1 U6545 ( .A1(n9446), .A2(n5457), .A3(n9445), .ZN(n12207) );
  NAND3_X1 U6546 ( .A1(n9412), .A2(n5457), .A3(n9411), .ZN(n12208) );
  NAND3_X1 U6547 ( .A1(n9305), .A2(n5457), .A3(n9304), .ZN(n12211) );
  NAND3_X1 U6548 ( .A1(n9374), .A2(n5457), .A3(n9373), .ZN(n12309) );
  NAND3_X1 U6549 ( .A1(n9240), .A2(n5457), .A3(n9239), .ZN(n12312) );
  NAND3_X1 U6550 ( .A1(n9272), .A2(n5457), .A3(n9271), .ZN(n12491) );
  NAND3_X1 U6551 ( .A1(net359513), .A2(net359680), .A3(net359515), .ZN(n12522)
         );
  INV_X4 U6552 ( .A(n6593), .ZN(n6597) );
  INV_X16 U6553 ( .A(n6598), .ZN(n6596) );
  OAI21_X2 U6554 ( .B1(n6562), .B2(n9516), .A(n6525), .ZN(n9520) );
  OAI21_X2 U6555 ( .B1(n6562), .B2(n9601), .A(n6527), .ZN(n9605) );
  INV_X4 U6556 ( .A(n13243), .ZN(n13246) );
  NAND3_X1 U6557 ( .A1(ifInst[30]), .A2(n13539), .A3(ifInst[28]), .ZN(n2054)
         );
  NOR2_X2 U6558 ( .A1(n13434), .A2(n13358), .ZN(n13360) );
  NOR2_X2 U6559 ( .A1(n6607), .A2(idOut_38_), .ZN(n3356) );
  INV_X16 U6560 ( .A(n6593), .ZN(n6594) );
  NAND3_X2 U6561 ( .A1(n13511), .A2(n13510), .A3(n13509), .ZN(n13512) );
  OAI21_X2 U6562 ( .B1(n6639), .B2(n6733), .A(n592), .ZN(n4183) );
  OAI21_X2 U6563 ( .B1(n6639), .B2(n6741), .A(n526), .ZN(n4185) );
  OAI21_X2 U6564 ( .B1(n6652), .B2(net367217), .A(n400), .ZN(n3930) );
  OAI21_X2 U6565 ( .B1(n6651), .B2(net367595), .A(n1103), .ZN(n3938) );
  OAI21_X2 U6566 ( .B1(n6651), .B2(n6708), .A(n835), .ZN(n3946) );
  OAI21_X2 U6567 ( .B1(n6652), .B2(n6741), .A(n534), .ZN(n3954) );
  OAI21_X2 U6568 ( .B1(n6638), .B2(n6711), .A(n793), .ZN(n4178) );
  NAND3_X2 U6569 ( .A1(n12949), .A2(n12948), .A3(n12947), .ZN(n4723) );
  NOR2_X2 U6570 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  OAI21_X2 U6571 ( .B1(n6649), .B2(n6679), .A(n1135), .ZN(n3961) );
  OAI21_X2 U6572 ( .B1(n6650), .B2(net367217), .A(n399), .ZN(n3963) );
  OAI21_X2 U6573 ( .B1(n6649), .B2(n6701), .A(n900), .ZN(n3977) );
  OAI21_X2 U6574 ( .B1(n6649), .B2(n6708), .A(n834), .ZN(n3979) );
  OAI21_X2 U6575 ( .B1(n6650), .B2(n6733), .A(n599), .ZN(n3985) );
  OAI21_X2 U6576 ( .B1(n6650), .B2(n6741), .A(n533), .ZN(n3987) );
  OAI21_X2 U6577 ( .B1(n5661), .B2(n6776), .A(n120), .ZN(n4167) );
  OAI21_X2 U6578 ( .B1(n6638), .B2(n6708), .A(n827), .ZN(n4177) );
  OAI21_X2 U6579 ( .B1(n6638), .B2(n6679), .A(n1128), .ZN(n4159) );
  OAI21_X2 U6580 ( .B1(n6638), .B2(n6701), .A(n893), .ZN(n4175) );
  OAI21_X2 U6581 ( .B1(n6638), .B2(n6705), .A(n860), .ZN(n4176) );
  NOR2_X2 U6582 ( .A1(n12224), .A2(net368481), .ZN(aluBoi_multBoi_N55) );
  NOR2_X2 U6583 ( .A1(n12331), .A2(net368481), .ZN(aluBoi_multBoi_N57) );
  NOR2_X2 U6584 ( .A1(n10067), .A2(n10066), .ZN(n10068) );
  NOR2_X2 U6585 ( .A1(n12222), .A2(net367631), .ZN(aluBoi_multBoi_N47) );
  NOR2_X2 U6586 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  OAI21_X2 U6587 ( .B1(n6628), .B2(n6698), .A(n922), .ZN(n4339) );
  OAI21_X2 U6588 ( .B1(n6636), .B2(n6699), .A(n926), .ZN(n4207) );
  OAI21_X2 U6589 ( .B1(n6624), .B2(n6705), .A(n853), .ZN(n4407) );
  OAI21_X2 U6590 ( .B1(n5655), .B2(n6757), .A(n331), .ZN(n4025) );
  OAI21_X2 U6591 ( .B1(n6655), .B2(n6713), .A(n770), .ZN(n3863) );
  OAI21_X2 U6592 ( .B1(n5651), .B2(n6758), .A(n301), .ZN(n3865) );
  OAI21_X2 U6593 ( .B1(n6667), .B2(n6749), .A(n411), .ZN(n3660) );
  OAI21_X2 U6594 ( .B1(n6625), .B2(n6733), .A(n585), .ZN(n4414) );
  OAI21_X2 U6595 ( .B1(n5682), .B2(n6684), .A(n1054), .ZN(n4434) );
  OAI21_X2 U6596 ( .B1(n6647), .B2(n6699), .A(n933), .ZN(n4009) );
  OAI21_X2 U6597 ( .B1(n6635), .B2(n6734), .A(n590), .ZN(n4249) );
  OAI21_X2 U6598 ( .B1(n6623), .B2(n6741), .A(n518), .ZN(n4449) );
  OAI21_X2 U6599 ( .B1(n6647), .B2(n6694), .A(n967), .ZN(n4008) );
  OAI21_X2 U6600 ( .B1(n6635), .B2(n6745), .A(n490), .ZN(n4252) );
  OAI21_X2 U6601 ( .B1(n6634), .B2(n6699), .A(n925), .ZN(n4240) );
  OAI21_X2 U6602 ( .B1(n6624), .B2(n6708), .A(n820), .ZN(n4408) );
  OAI21_X2 U6603 ( .B1(n6664), .B2(n6697), .A(n912), .ZN(n3679) );
  OAI21_X2 U6604 ( .B1(n5652), .B2(n6756), .A(n334), .ZN(n3926) );
  OAI21_X2 U6605 ( .B1(n6623), .B2(n6753), .A(n351), .ZN(n4453) );
  OAI21_X2 U6606 ( .B1(n6620), .B2(net367215), .A(n381), .ZN(n4491) );
  OAI21_X2 U6607 ( .B1(n6675), .B2(n6751), .A(n427), .ZN(n3528) );
  OAI21_X2 U6608 ( .B1(n6675), .B2(n439), .A(n460), .ZN(n3527) );
  OAI21_X2 U6609 ( .B1(n5659), .B2(n6774), .A(n156), .ZN(n3506) );
  OAI21_X2 U6610 ( .B1(n5673), .B2(n6772), .A(n138), .ZN(n3704) );
  OAI21_X2 U6611 ( .B1(n6675), .B2(n340), .A(n361), .ZN(n3529) );
  OAI21_X2 U6612 ( .B1(n6779), .B2(n5688), .A(n46), .ZN(n3607) );
  OAI21_X2 U6613 ( .B1(n6660), .B2(n6697), .A(n910), .ZN(n3745) );
  OAI21_X2 U6614 ( .B1(n6668), .B2(net367593), .A(n1082), .ZN(n3608) );
  OAI21_X2 U6615 ( .B1(n6668), .B2(n6686), .A(n1015), .ZN(n3610) );
  OAI21_X2 U6616 ( .B1(n5674), .B2(n6755), .A(n308), .ZN(n3761) );
  OAI21_X2 U6617 ( .B1(n6662), .B2(n6689), .A(n978), .ZN(n3710) );
  OAI21_X2 U6618 ( .B1(n6662), .B2(n6683), .A(n1046), .ZN(n3708) );
  OAI21_X2 U6619 ( .B1(n6662), .B2(n6693), .A(n945), .ZN(n3711) );
  OAI21_X2 U6620 ( .B1(n5688), .B2(n6768), .A(n176), .ZN(n3604) );
  OAI21_X2 U6621 ( .B1(n6669), .B2(n6717), .A(n714), .ZN(n3618) );
  OAI21_X2 U6622 ( .B1(n5659), .B2(n6757), .A(n327), .ZN(n3530) );
  OAI21_X2 U6623 ( .B1(n5669), .B2(n6756), .A(n316), .ZN(n3563) );
  OAI21_X2 U6624 ( .B1(n6668), .B2(n6689), .A(n981), .ZN(n3611) );
  OAI21_X2 U6625 ( .B1(n6659), .B2(n6717), .A(n709), .ZN(n3783) );
  OAI21_X2 U6626 ( .B1(n6635), .B2(n6740), .A(n524), .ZN(n4251) );
  OAI21_X2 U6627 ( .B1(n6634), .B2(n6709), .A(n825), .ZN(n4243) );
  OAI21_X2 U6628 ( .B1(n6627), .B2(n6733), .A(n586), .ZN(n4381) );
  OAI21_X2 U6629 ( .B1(n6626), .B2(n6701), .A(n887), .ZN(n4373) );
  OAI21_X2 U6630 ( .B1(n6654), .B2(n6747), .A(n467), .ZN(n3923) );
  OAI21_X2 U6631 ( .B1(n6654), .B2(n6753), .A(n368), .ZN(n3925) );
  OAI21_X2 U6632 ( .B1(n6635), .B2(n6730), .A(n625), .ZN(n4248) );
  OAI21_X2 U6633 ( .B1(n5663), .B2(n6757), .A(n323), .ZN(n4256) );
  OAI21_X2 U6634 ( .B1(n6635), .B2(n6753), .A(n357), .ZN(n4255) );
  OAI21_X2 U6635 ( .B1(n6635), .B2(n6727), .A(n659), .ZN(n4247) );
  OAI21_X2 U6636 ( .B1(n6625), .B2(n6741), .A(n519), .ZN(n4416) );
  OAI21_X2 U6637 ( .B1(n6624), .B2(net367595), .A(n1088), .ZN(n4400) );
  OAI21_X2 U6638 ( .B1(n6658), .B2(n6736), .A(n571), .ZN(n3821) );
  OAI21_X2 U6639 ( .B1(n6658), .B2(n6710), .A(n805), .ZN(n3815) );
  OAI21_X2 U6640 ( .B1(n6658), .B2(n6693), .A(n973), .ZN(n3810) );
  OAI21_X2 U6641 ( .B1(n6658), .B2(n6722), .A(n706), .ZN(n3817) );
  OAI21_X2 U6642 ( .B1(n6658), .B2(n6740), .A(n538), .ZN(n3822) );
  OAI21_X2 U6643 ( .B1(n6658), .B2(n6683), .A(n1074), .ZN(n3807) );
  OAI21_X2 U6644 ( .B1(n5649), .B2(n6758), .A(n303), .ZN(n3799) );
  OAI21_X2 U6645 ( .B1(n5675), .B2(n6772), .A(n136), .ZN(n3770) );
  OAI21_X2 U6646 ( .B1(n6779), .B2(n5675), .A(n36), .ZN(n3772) );
  OAI21_X2 U6647 ( .B1(n6659), .B2(n6689), .A(n976), .ZN(n3776) );
  OAI21_X2 U6648 ( .B1(n6669), .B2(n6736), .A(n546), .ZN(n3623) );
  OAI21_X2 U6649 ( .B1(n6668), .B2(n6693), .A(n948), .ZN(n3612) );
  OAI21_X2 U6650 ( .B1(n6659), .B2(n6693), .A(n943), .ZN(n3777) );
  OAI21_X2 U6651 ( .B1(n6669), .B2(n6740), .A(n513), .ZN(n3624) );
  OAI21_X2 U6652 ( .B1(n5688), .B2(n6772), .A(n141), .ZN(n3605) );
  OAI21_X2 U6653 ( .B1(n6668), .B2(n6683), .A(n1049), .ZN(n3609) );
  OAI21_X2 U6654 ( .B1(n6659), .B2(n6740), .A(n508), .ZN(n3789) );
  OAI21_X2 U6655 ( .B1(n6658), .B2(n6728), .A(n639), .ZN(n3819) );
  OAI21_X2 U6656 ( .B1(n6658), .B2(n6743), .A(n504), .ZN(n3823) );
  OAI21_X2 U6657 ( .B1(n6662), .B2(n6697), .A(n911), .ZN(n3712) );
  OAI21_X2 U6658 ( .B1(n6658), .B2(n6749), .A(n437), .ZN(n3825) );
  OAI21_X2 U6659 ( .B1(n6658), .B2(n6697), .A(n939), .ZN(n3811) );
  OAI21_X2 U6660 ( .B1(n6670), .B2(n6697), .A(n915), .ZN(n3580) );
  OAI21_X2 U6661 ( .B1(n6670), .B2(n6693), .A(n949), .ZN(n3579) );
  OAI21_X2 U6662 ( .B1(n6671), .B2(n6743), .A(n480), .ZN(n3592) );
  OAI21_X2 U6663 ( .B1(n6671), .B2(n6749), .A(n413), .ZN(n3594) );
  OAI21_X2 U6664 ( .B1(n6671), .B2(n6752), .A(n347), .ZN(n3595) );
  OAI21_X2 U6665 ( .B1(n6659), .B2(n6697), .A(n909), .ZN(n3778) );
  OAI21_X2 U6666 ( .B1(n5675), .B2(n6749), .A(n407), .ZN(n3792) );
  OAI21_X2 U6667 ( .B1(n6668), .B2(n6697), .A(n914), .ZN(n3613) );
  OAI21_X2 U6668 ( .B1(n5649), .B2(n6755), .A(n337), .ZN(n3827) );
  OAI21_X2 U6669 ( .B1(n5649), .B2(n6752), .A(n371), .ZN(n3826) );
  OAI21_X2 U6670 ( .B1(n6659), .B2(n6752), .A(n341), .ZN(n3793) );
  OAI21_X2 U6671 ( .B1(n6659), .B2(n6725), .A(n643), .ZN(n3785) );
  OAI21_X2 U6672 ( .B1(n6669), .B2(n6752), .A(n346), .ZN(n3628) );
  OAI21_X2 U6673 ( .B1(n6669), .B2(n6725), .A(n648), .ZN(n3620) );
  OAI21_X2 U6674 ( .B1(n6659), .B2(n6743), .A(n474), .ZN(n3790) );
  OAI21_X2 U6675 ( .B1(n6659), .B2(n6710), .A(n775), .ZN(n3782) );
  OAI21_X2 U6676 ( .B1(n5688), .B2(n6755), .A(n312), .ZN(n3629) );
  OAI21_X2 U6677 ( .B1(n6669), .B2(n6728), .A(n614), .ZN(n3621) );
  OAI21_X2 U6678 ( .B1(n6669), .B2(n6743), .A(n479), .ZN(n3625) );
  OAI21_X2 U6679 ( .B1(n6668), .B2(n6710), .A(n780), .ZN(n3617) );
  OAI21_X2 U6680 ( .B1(n5671), .B2(n6755), .A(n313), .ZN(n3596) );
  OAI21_X2 U6681 ( .B1(n6671), .B2(n6728), .A(n615), .ZN(n3588) );
  OAI21_X2 U6682 ( .B1(n5675), .B2(n6755), .A(n307), .ZN(n3794) );
  OAI21_X2 U6683 ( .B1(n6659), .B2(n6728), .A(n609), .ZN(n3786) );
  OAI21_X2 U6684 ( .B1(n6669), .B2(n6749), .A(n412), .ZN(n3627) );
  OAI21_X2 U6685 ( .B1(n6669), .B2(n6722), .A(n681), .ZN(n3619) );
  NOR2_X2 U6686 ( .A1(n10094), .A2(n10093), .ZN(n10095) );
  NAND3_X2 U6687 ( .A1(n10133), .A2(n10132), .A3(n10131), .ZN(n4603) );
  AOI21_X2 U6688 ( .B1(iaddr[9]), .B2(n10301), .A(n10300), .ZN(n10302) );
  AOI21_X1 U6689 ( .B1(n6571), .B2(n12883), .A(n6434), .ZN(n10365) );
  NAND3_X2 U6690 ( .A1(n10411), .A2(n10410), .A3(n10409), .ZN(n4713) );
  AOI21_X2 U6691 ( .B1(n6576), .B2(n10405), .A(n10404), .ZN(n10411) );
  OAI21_X2 U6692 ( .B1(net100619), .B2(n5691), .A(n2105), .ZN(n4873) );
  OAI21_X2 U6693 ( .B1(idOut_20_), .B2(n2840), .A(n2841), .ZN(
        aluBoi_condBoi_N25) );
  NAND3_X2 U6694 ( .A1(n2842), .A2(n5715), .A3(n13575), .ZN(n2841) );
  NOR2_X1 U6695 ( .A1(net368481), .A2(n5471), .ZN(aluBoi_multBoi_N6) );
  NOR2_X2 U6696 ( .A1(n10679), .A2(n10678), .ZN(n10681) );
  NOR2_X2 U6697 ( .A1(net367631), .A2(n12321), .ZN(aluBoi_multBoi_N41) );
  NOR3_X2 U6698 ( .A1(n12497), .A2(net368481), .A3(n12496), .ZN(
        aluBoi_multBoi_N40) );
  NOR2_X1 U6699 ( .A1(n12494), .A2(n12493), .ZN(n12497) );
  NOR2_X2 U6700 ( .A1(aluBoi_multBoi_count_0_), .A2(aluBoi_multBoi_count_1_), 
        .ZN(n2203) );
  OAI21_X2 U6701 ( .B1(n6676), .B2(n6678), .A(n1141), .ZN(n3466) );
  OAI21_X2 U6702 ( .B1(n6676), .B2(n6713), .A(n773), .ZN(n3467) );
  OAI21_X2 U6703 ( .B1(n6677), .B2(net367215), .A(n405), .ZN(n3468) );
  OAI21_X2 U6704 ( .B1(n6677), .B2(n6758), .A(n304), .ZN(n3469) );
  OAI21_X2 U6705 ( .B1(n5648), .B2(n6761), .A(n269), .ZN(n3470) );
  OAI21_X2 U6706 ( .B1(n6676), .B2(n6765), .A(n236), .ZN(n3471) );
  OAI21_X2 U6707 ( .B1(n5648), .B2(n6768), .A(n202), .ZN(n3472) );
  OAI21_X2 U6708 ( .B1(n5648), .B2(n6772), .A(n167), .ZN(n3473) );
  OAI21_X2 U6709 ( .B1(n5648), .B2(n6775), .A(n133), .ZN(n3474) );
  OAI21_X2 U6710 ( .B1(n6779), .B2(n5648), .A(n98), .ZN(n3475) );
  OAI21_X2 U6711 ( .B1(n6676), .B2(net367593), .A(n1108), .ZN(n3476) );
  OAI21_X2 U6712 ( .B1(n6676), .B2(n6683), .A(n1075), .ZN(n3477) );
  OAI21_X2 U6713 ( .B1(n6676), .B2(n6686), .A(n1041), .ZN(n3478) );
  OAI21_X2 U6714 ( .B1(n6676), .B2(n6689), .A(n1007), .ZN(n3479) );
  OAI21_X2 U6715 ( .B1(n6676), .B2(n6693), .A(n974), .ZN(n3480) );
  OAI21_X2 U6716 ( .B1(n6676), .B2(n6697), .A(n940), .ZN(n3481) );
  OAI21_X2 U6717 ( .B1(n6676), .B2(n6700), .A(n906), .ZN(n3482) );
  OAI21_X2 U6718 ( .B1(n6676), .B2(n6704), .A(n873), .ZN(n3483) );
  OAI21_X2 U6719 ( .B1(n6676), .B2(n6707), .A(n840), .ZN(n3484) );
  OAI21_X2 U6720 ( .B1(n6676), .B2(n6710), .A(n806), .ZN(n3485) );
  OAI21_X2 U6721 ( .B1(n6677), .B2(n6717), .A(n740), .ZN(n3486) );
  OAI21_X2 U6722 ( .B1(n6677), .B2(n6722), .A(n707), .ZN(n3487) );
  OAI21_X2 U6723 ( .B1(n6677), .B2(n6725), .A(n674), .ZN(n3488) );
  OAI21_X2 U6724 ( .B1(n6677), .B2(n6728), .A(n640), .ZN(n3489) );
  OAI21_X2 U6725 ( .B1(n6677), .B2(n6732), .A(n605), .ZN(n3490) );
  OAI21_X2 U6726 ( .B1(n6677), .B2(n6736), .A(n572), .ZN(n3491) );
  OAI21_X2 U6727 ( .B1(n6677), .B2(n6740), .A(n539), .ZN(n3492) );
  OAI21_X2 U6728 ( .B1(n6677), .B2(n6743), .A(n505), .ZN(n3493) );
  OAI21_X2 U6729 ( .B1(n6677), .B2(n439), .A(n471), .ZN(n3494) );
  OAI21_X2 U6730 ( .B1(n6677), .B2(n6749), .A(n438), .ZN(n3495) );
  OAI21_X2 U6731 ( .B1(n6677), .B2(n6752), .A(n372), .ZN(n3496) );
  OAI21_X2 U6732 ( .B1(n6676), .B2(n6755), .A(n338), .ZN(n3497) );
  AOI21_X2 U6733 ( .B1(drData[31]), .B2(n1158), .A(n13673), .ZN(n1157) );
  OAI21_X2 U6734 ( .B1(n6674), .B2(n6678), .A(n1130), .ZN(n3499) );
  OAI21_X2 U6735 ( .B1(n6674), .B2(n6713), .A(n762), .ZN(n3500) );
  OAI21_X2 U6736 ( .B1(n6675), .B2(n373), .A(n394), .ZN(n3501) );
  OAI21_X2 U6737 ( .B1(n6674), .B2(n6760), .A(n293), .ZN(n3502) );
  OAI21_X2 U6738 ( .B1(n6674), .B2(n237), .A(n258), .ZN(n3503) );
  OAI21_X2 U6739 ( .B1(n6675), .B2(n6767), .A(n225), .ZN(n3504) );
  OAI21_X2 U6740 ( .B1(n5659), .B2(n6770), .A(n191), .ZN(n3505) );
  OAI21_X2 U6741 ( .B1(n5659), .B2(n6777), .A(n122), .ZN(n3507) );
  OAI21_X2 U6742 ( .B1(n6780), .B2(n5659), .A(n76), .ZN(n3508) );
  OAI21_X2 U6743 ( .B1(n6674), .B2(net367597), .A(n1097), .ZN(n3509) );
  OAI21_X2 U6744 ( .B1(n6674), .B2(n6684), .A(n1064), .ZN(n3510) );
  OAI21_X2 U6745 ( .B1(n6674), .B2(n6688), .A(n1030), .ZN(n3511) );
  OAI21_X2 U6746 ( .B1(n6674), .B2(n6691), .A(n996), .ZN(n3512) );
  OAI21_X2 U6747 ( .B1(n6674), .B2(n942), .A(n963), .ZN(n3513) );
  OAI21_X2 U6748 ( .B1(n6674), .B2(n6699), .A(n929), .ZN(n3514) );
  OAI21_X2 U6749 ( .B1(n6674), .B2(n6702), .A(n895), .ZN(n3515) );
  OAI21_X2 U6750 ( .B1(n6674), .B2(n6706), .A(n862), .ZN(n3516) );
  OAI21_X2 U6751 ( .B1(n6674), .B2(n6709), .A(n829), .ZN(n3517) );
  OAI21_X2 U6752 ( .B1(n6674), .B2(n6712), .A(n795), .ZN(n3518) );
  OAI21_X2 U6753 ( .B1(n6675), .B2(n708), .A(n729), .ZN(n3519) );
  OAI21_X2 U6754 ( .B1(n6675), .B2(n675), .A(n696), .ZN(n3520) );
  OAI21_X2 U6755 ( .B1(n6675), .B2(n6727), .A(n663), .ZN(n3521) );
  OAI21_X2 U6756 ( .B1(n6675), .B2(n6730), .A(n629), .ZN(n3522) );
  OAI21_X2 U6757 ( .B1(n6675), .B2(n6734), .A(n594), .ZN(n3523) );
  OAI21_X2 U6758 ( .B1(n6675), .B2(n540), .A(n561), .ZN(n3524) );
  OAI21_X2 U6759 ( .B1(n6675), .B2(n507), .A(n528), .ZN(n3525) );
  OAI21_X2 U6760 ( .B1(n6675), .B2(n6745), .A(n494), .ZN(n3526) );
  AOI21_X2 U6761 ( .B1(drData[30]), .B2(n1158), .A(n13673), .ZN(n1162) );
  OAI21_X2 U6762 ( .B1(n6672), .B2(n6679), .A(n1119), .ZN(n3532) );
  OAI21_X2 U6763 ( .B1(n6672), .B2(n6714), .A(n751), .ZN(n3533) );
  OAI21_X2 U6764 ( .B1(n6673), .B2(net367217), .A(n383), .ZN(n3534) );
  OAI21_X2 U6765 ( .B1(n6672), .B2(n6759), .A(n282), .ZN(n3535) );
  OAI21_X2 U6766 ( .B1(n5669), .B2(n6762), .A(n247), .ZN(n3536) );
  OAI21_X2 U6767 ( .B1(n6673), .B2(n6766), .A(n214), .ZN(n3537) );
  OAI21_X2 U6768 ( .B1(n5669), .B2(n6769), .A(n180), .ZN(n3538) );
  OAI21_X2 U6769 ( .B1(n6672), .B2(n6773), .A(n145), .ZN(n3539) );
  OAI21_X2 U6770 ( .B1(n5669), .B2(n6776), .A(n111), .ZN(n3540) );
  OAI21_X2 U6771 ( .B1(n6780), .B2(n5669), .A(n54), .ZN(n3541) );
  OAI21_X2 U6772 ( .B1(n6672), .B2(net367595), .A(n1086), .ZN(n3542) );
  OAI21_X2 U6773 ( .B1(n6672), .B2(n6684), .A(n1053), .ZN(n3543) );
  OAI21_X2 U6774 ( .B1(n6672), .B2(n6687), .A(n1019), .ZN(n3544) );
  OAI21_X2 U6775 ( .B1(n6672), .B2(n6690), .A(n985), .ZN(n3545) );
  OAI21_X2 U6776 ( .B1(n6672), .B2(n6694), .A(n952), .ZN(n3546) );
  OAI21_X2 U6777 ( .B1(n6672), .B2(n6698), .A(n918), .ZN(n3547) );
  OAI21_X2 U6778 ( .B1(n6672), .B2(n6701), .A(n884), .ZN(n3548) );
  OAI21_X2 U6779 ( .B1(n6672), .B2(n6705), .A(n851), .ZN(n3549) );
  OAI21_X2 U6780 ( .B1(n6672), .B2(n6708), .A(n818), .ZN(n3550) );
  OAI21_X2 U6781 ( .B1(n6672), .B2(n6711), .A(n784), .ZN(n3551) );
  OAI21_X2 U6782 ( .B1(n6673), .B2(n6718), .A(n718), .ZN(n3552) );
  OAI21_X2 U6783 ( .B1(n6673), .B2(n6723), .A(n685), .ZN(n3553) );
  OAI21_X2 U6784 ( .B1(n6673), .B2(n6726), .A(n652), .ZN(n3554) );
  OAI21_X2 U6785 ( .B1(n6673), .B2(n6729), .A(n618), .ZN(n3555) );
  OAI21_X2 U6786 ( .B1(n6673), .B2(n6733), .A(n583), .ZN(n3556) );
  OAI21_X2 U6787 ( .B1(n6673), .B2(n6737), .A(n550), .ZN(n3557) );
  OAI21_X2 U6788 ( .B1(n6673), .B2(n6741), .A(n517), .ZN(n3558) );
  OAI21_X2 U6789 ( .B1(n6673), .B2(n6744), .A(n483), .ZN(n3559) );
  OAI21_X2 U6790 ( .B1(n6673), .B2(n6747), .A(n449), .ZN(n3560) );
  OAI21_X2 U6791 ( .B1(n6673), .B2(n6750), .A(n416), .ZN(n3561) );
  OAI21_X2 U6792 ( .B1(n6673), .B2(n6753), .A(n350), .ZN(n3562) );
  AOI21_X2 U6793 ( .B1(drData[29]), .B2(n1158), .A(n13673), .ZN(n1165) );
  OAI21_X2 U6794 ( .B1(n6670), .B2(n6678), .A(n1116), .ZN(n3565) );
  OAI21_X2 U6795 ( .B1(n6670), .B2(n6713), .A(n748), .ZN(n3566) );
  OAI21_X2 U6796 ( .B1(n6671), .B2(net367215), .A(n380), .ZN(n3567) );
  OAI21_X2 U6797 ( .B1(n6670), .B2(n6758), .A(n279), .ZN(n3568) );
  OAI21_X2 U6798 ( .B1(n5671), .B2(n6761), .A(n244), .ZN(n3569) );
  OAI21_X2 U6799 ( .B1(n6671), .B2(n6765), .A(n211), .ZN(n3570) );
  OAI21_X2 U6800 ( .B1(n5671), .B2(n6768), .A(n177), .ZN(n3571) );
  OAI21_X2 U6801 ( .B1(n6670), .B2(n6772), .A(n142), .ZN(n3572) );
  OAI21_X2 U6802 ( .B1(n5671), .B2(n6775), .A(n108), .ZN(n3573) );
  OAI21_X2 U6803 ( .B1(n6779), .B2(n5671), .A(n48), .ZN(n3574) );
  OAI21_X2 U6804 ( .B1(n6670), .B2(net367593), .A(n1083), .ZN(n3575) );
  OAI21_X2 U6805 ( .B1(n6670), .B2(n6683), .A(n1050), .ZN(n3576) );
  OAI21_X2 U6806 ( .B1(n6670), .B2(n6686), .A(n1016), .ZN(n3577) );
  OAI21_X2 U6807 ( .B1(n6670), .B2(n6689), .A(n982), .ZN(n3578) );
  OAI21_X2 U6808 ( .B1(n6670), .B2(n6700), .A(n881), .ZN(n3581) );
  OAI21_X2 U6809 ( .B1(n6670), .B2(n6704), .A(n848), .ZN(n3582) );
  OAI21_X2 U6810 ( .B1(n6670), .B2(n6707), .A(n815), .ZN(n3583) );
  OAI21_X2 U6811 ( .B1(n6670), .B2(n6710), .A(n781), .ZN(n3584) );
  OAI21_X2 U6812 ( .B1(n6671), .B2(n6717), .A(n715), .ZN(n3585) );
  OAI21_X2 U6813 ( .B1(n6671), .B2(n6722), .A(n682), .ZN(n3586) );
  OAI21_X2 U6814 ( .B1(n6671), .B2(n6725), .A(n649), .ZN(n3587) );
  OAI21_X2 U6815 ( .B1(n6671), .B2(n6732), .A(n580), .ZN(n3589) );
  OAI21_X2 U6816 ( .B1(n6671), .B2(n6736), .A(n547), .ZN(n3590) );
  OAI21_X2 U6817 ( .B1(n6671), .B2(n6740), .A(n514), .ZN(n3591) );
  OAI21_X2 U6818 ( .B1(n6671), .B2(n439), .A(n446), .ZN(n3593) );
  AOI21_X2 U6819 ( .B1(drData[28]), .B2(n1158), .A(n13673), .ZN(n1168) );
  OAI21_X2 U6820 ( .B1(n6668), .B2(n6678), .A(n1115), .ZN(n3598) );
  OAI21_X2 U6821 ( .B1(n6668), .B2(n6713), .A(n747), .ZN(n3599) );
  OAI21_X2 U6822 ( .B1(n6669), .B2(net367215), .A(n379), .ZN(n3600) );
  OAI21_X2 U6823 ( .B1(n6669), .B2(n6761), .A(n243), .ZN(n3602) );
  OAI21_X2 U6824 ( .B1(n6668), .B2(n6775), .A(n107), .ZN(n3606) );
  OAI21_X2 U6825 ( .B1(n6668), .B2(n6700), .A(n880), .ZN(n3614) );
  OAI21_X2 U6826 ( .B1(n6668), .B2(n6707), .A(n814), .ZN(n3616) );
  OAI21_X2 U6827 ( .B1(n6669), .B2(n6732), .A(n579), .ZN(n3622) );
  AOI21_X2 U6828 ( .B1(drData[27]), .B2(n1158), .A(n13673), .ZN(n1171) );
  OAI21_X2 U6829 ( .B1(n6666), .B2(n6678), .A(n1114), .ZN(n3631) );
  OAI21_X2 U6830 ( .B1(n6666), .B2(n6713), .A(n746), .ZN(n3632) );
  OAI21_X2 U6831 ( .B1(n6667), .B2(net367215), .A(n378), .ZN(n3633) );
  OAI21_X2 U6832 ( .B1(n6666), .B2(n6758), .A(n277), .ZN(n3634) );
  OAI21_X2 U6833 ( .B1(n5672), .B2(n6761), .A(n242), .ZN(n3635) );
  OAI21_X2 U6834 ( .B1(n6667), .B2(n6765), .A(n209), .ZN(n3636) );
  OAI21_X2 U6835 ( .B1(n5672), .B2(n6768), .A(n175), .ZN(n3637) );
  OAI21_X2 U6836 ( .B1(n6666), .B2(n6772), .A(n140), .ZN(n3638) );
  OAI21_X2 U6837 ( .B1(n5672), .B2(n6775), .A(n106), .ZN(n3639) );
  OAI21_X2 U6838 ( .B1(n6779), .B2(n5672), .A(n44), .ZN(n3640) );
  OAI21_X2 U6839 ( .B1(n6666), .B2(net367593), .A(n1081), .ZN(n3641) );
  OAI21_X2 U6840 ( .B1(n6666), .B2(n6683), .A(n1048), .ZN(n3642) );
  OAI21_X2 U6841 ( .B1(n6666), .B2(n6686), .A(n1014), .ZN(n3643) );
  OAI21_X2 U6842 ( .B1(n6666), .B2(n6689), .A(n980), .ZN(n3644) );
  OAI21_X2 U6843 ( .B1(n6666), .B2(n6693), .A(n947), .ZN(n3645) );
  OAI21_X2 U6844 ( .B1(n6666), .B2(n6697), .A(n913), .ZN(n3646) );
  OAI21_X2 U6845 ( .B1(n6666), .B2(n6700), .A(n879), .ZN(n3647) );
  OAI21_X2 U6846 ( .B1(n6666), .B2(n6704), .A(n846), .ZN(n3648) );
  OAI21_X2 U6847 ( .B1(n6666), .B2(n6707), .A(n813), .ZN(n3649) );
  OAI21_X2 U6848 ( .B1(n6666), .B2(n6710), .A(n779), .ZN(n3650) );
  OAI21_X2 U6849 ( .B1(n6667), .B2(n6717), .A(n713), .ZN(n3651) );
  OAI21_X2 U6850 ( .B1(n6667), .B2(n6722), .A(n680), .ZN(n3652) );
  OAI21_X2 U6851 ( .B1(n6667), .B2(n6725), .A(n647), .ZN(n3653) );
  OAI21_X2 U6852 ( .B1(n6667), .B2(n6728), .A(n613), .ZN(n3654) );
  OAI21_X2 U6853 ( .B1(n6667), .B2(n6732), .A(n578), .ZN(n3655) );
  OAI21_X2 U6854 ( .B1(n6667), .B2(n6736), .A(n545), .ZN(n3656) );
  OAI21_X2 U6855 ( .B1(n6667), .B2(n6740), .A(n512), .ZN(n3657) );
  OAI21_X2 U6856 ( .B1(n6667), .B2(n6743), .A(n478), .ZN(n3658) );
  OAI21_X2 U6857 ( .B1(n6667), .B2(n439), .A(n444), .ZN(n3659) );
  OAI21_X2 U6858 ( .B1(n6667), .B2(n6752), .A(n345), .ZN(n3661) );
  OAI21_X2 U6859 ( .B1(n5672), .B2(n6755), .A(n311), .ZN(n3662) );
  AOI21_X2 U6860 ( .B1(drData[26]), .B2(n1158), .A(n13673), .ZN(n1174) );
  OAI21_X2 U6861 ( .B1(n6664), .B2(n6678), .A(n1113), .ZN(n3664) );
  OAI21_X2 U6862 ( .B1(n6664), .B2(n6713), .A(n745), .ZN(n3665) );
  OAI21_X2 U6863 ( .B1(n6665), .B2(net367215), .A(n377), .ZN(n3666) );
  OAI21_X2 U6864 ( .B1(n6665), .B2(n6758), .A(n276), .ZN(n3667) );
  OAI21_X2 U6865 ( .B1(n5684), .B2(n6761), .A(n241), .ZN(n3668) );
  OAI21_X2 U6866 ( .B1(n6664), .B2(n6765), .A(n208), .ZN(n3669) );
  OAI21_X2 U6867 ( .B1(n5684), .B2(n6768), .A(n174), .ZN(n3670) );
  OAI21_X2 U6868 ( .B1(n6665), .B2(n6772), .A(n139), .ZN(n3671) );
  OAI21_X2 U6869 ( .B1(n5684), .B2(n6775), .A(n105), .ZN(n3672) );
  OAI21_X2 U6870 ( .B1(n6779), .B2(n5684), .A(n42), .ZN(n3673) );
  OAI21_X2 U6871 ( .B1(n6664), .B2(net367593), .A(n1080), .ZN(n3674) );
  OAI21_X2 U6872 ( .B1(n6664), .B2(n6683), .A(n1047), .ZN(n3675) );
  OAI21_X2 U6873 ( .B1(n6664), .B2(n6686), .A(n1013), .ZN(n3676) );
  OAI21_X2 U6874 ( .B1(n6664), .B2(n6689), .A(n979), .ZN(n3677) );
  OAI21_X2 U6875 ( .B1(n6664), .B2(n6693), .A(n946), .ZN(n3678) );
  OAI21_X2 U6876 ( .B1(n6664), .B2(n6700), .A(n878), .ZN(n3680) );
  OAI21_X2 U6877 ( .B1(n6664), .B2(n6704), .A(n845), .ZN(n3681) );
  OAI21_X2 U6878 ( .B1(n6664), .B2(n6707), .A(n812), .ZN(n3682) );
  OAI21_X2 U6879 ( .B1(n6664), .B2(n6710), .A(n778), .ZN(n3683) );
  OAI21_X2 U6880 ( .B1(n6665), .B2(n6717), .A(n712), .ZN(n3684) );
  OAI21_X2 U6881 ( .B1(n6665), .B2(n6722), .A(n679), .ZN(n3685) );
  OAI21_X2 U6882 ( .B1(n6665), .B2(n6725), .A(n646), .ZN(n3686) );
  OAI21_X2 U6883 ( .B1(n6665), .B2(n6728), .A(n612), .ZN(n3687) );
  OAI21_X2 U6884 ( .B1(n6665), .B2(n6732), .A(n577), .ZN(n3688) );
  OAI21_X2 U6885 ( .B1(n6665), .B2(n6736), .A(n544), .ZN(n3689) );
  OAI21_X2 U6886 ( .B1(n6665), .B2(n6740), .A(n511), .ZN(n3690) );
  OAI21_X2 U6887 ( .B1(n6665), .B2(n6743), .A(n477), .ZN(n3691) );
  OAI21_X2 U6888 ( .B1(n6665), .B2(n439), .A(n443), .ZN(n3692) );
  OAI21_X2 U6889 ( .B1(n6665), .B2(n6749), .A(n410), .ZN(n3693) );
  OAI21_X2 U6890 ( .B1(n6665), .B2(n6752), .A(n344), .ZN(n3694) );
  AOI21_X2 U6891 ( .B1(drData[25]), .B2(n1158), .A(n13673), .ZN(n1177) );
  OAI21_X2 U6892 ( .B1(n6662), .B2(n6678), .A(n1112), .ZN(n3697) );
  OAI21_X2 U6893 ( .B1(n6662), .B2(n6713), .A(n744), .ZN(n3698) );
  OAI21_X2 U6894 ( .B1(n6663), .B2(net367215), .A(n376), .ZN(n3699) );
  OAI21_X2 U6895 ( .B1(n6662), .B2(n6758), .A(n275), .ZN(n3700) );
  OAI21_X2 U6896 ( .B1(n5673), .B2(n6761), .A(n240), .ZN(n3701) );
  OAI21_X2 U6897 ( .B1(n6663), .B2(n6765), .A(n207), .ZN(n3702) );
  OAI21_X2 U6898 ( .B1(n5673), .B2(n6768), .A(n173), .ZN(n3703) );
  OAI21_X2 U6899 ( .B1(n5673), .B2(n6775), .A(n104), .ZN(n3705) );
  OAI21_X2 U6900 ( .B1(n6779), .B2(n5673), .A(n40), .ZN(n3706) );
  OAI21_X2 U6901 ( .B1(n6662), .B2(net367593), .A(n1079), .ZN(n3707) );
  OAI21_X2 U6902 ( .B1(n6662), .B2(n6686), .A(n1012), .ZN(n3709) );
  OAI21_X2 U6903 ( .B1(n6662), .B2(n6700), .A(n877), .ZN(n3713) );
  OAI21_X2 U6904 ( .B1(n6662), .B2(n6704), .A(n844), .ZN(n3714) );
  OAI21_X2 U6905 ( .B1(n6662), .B2(n6707), .A(n811), .ZN(n3715) );
  OAI21_X2 U6906 ( .B1(n6662), .B2(n6710), .A(n777), .ZN(n3716) );
  OAI21_X2 U6907 ( .B1(n6663), .B2(n6717), .A(n711), .ZN(n3717) );
  OAI21_X2 U6908 ( .B1(n6663), .B2(n6722), .A(n678), .ZN(n3718) );
  OAI21_X2 U6909 ( .B1(n6663), .B2(n6725), .A(n645), .ZN(n3719) );
  OAI21_X2 U6910 ( .B1(n6663), .B2(n6728), .A(n611), .ZN(n3720) );
  OAI21_X2 U6911 ( .B1(n6663), .B2(n6732), .A(n576), .ZN(n3721) );
  OAI21_X2 U6912 ( .B1(n6663), .B2(n6736), .A(n543), .ZN(n3722) );
  OAI21_X2 U6913 ( .B1(n6663), .B2(n6740), .A(n510), .ZN(n3723) );
  OAI21_X2 U6914 ( .B1(n6663), .B2(n6743), .A(n476), .ZN(n3724) );
  OAI21_X2 U6915 ( .B1(n6663), .B2(n439), .A(n442), .ZN(n3725) );
  OAI21_X2 U6916 ( .B1(n6663), .B2(n6749), .A(n409), .ZN(n3726) );
  OAI21_X2 U6917 ( .B1(n6663), .B2(n6752), .A(n343), .ZN(n3727) );
  OAI21_X2 U6918 ( .B1(n6663), .B2(n6755), .A(n309), .ZN(n3728) );
  AOI21_X2 U6919 ( .B1(drData[24]), .B2(n1158), .A(n13673), .ZN(n1180) );
  OAI21_X2 U6920 ( .B1(n6660), .B2(n6678), .A(n1111), .ZN(n3730) );
  OAI21_X2 U6921 ( .B1(n6660), .B2(n6713), .A(n743), .ZN(n3731) );
  OAI21_X2 U6922 ( .B1(n6661), .B2(net367215), .A(n375), .ZN(n3732) );
  OAI21_X2 U6923 ( .B1(n6661), .B2(n6758), .A(n274), .ZN(n3733) );
  OAI21_X2 U6924 ( .B1(n5674), .B2(n6761), .A(n239), .ZN(n3734) );
  OAI21_X2 U6925 ( .B1(n6660), .B2(n6765), .A(n206), .ZN(n3735) );
  OAI21_X2 U6926 ( .B1(n5674), .B2(n6768), .A(n172), .ZN(n3736) );
  OAI21_X2 U6927 ( .B1(n6661), .B2(n6772), .A(n137), .ZN(n3737) );
  OAI21_X2 U6928 ( .B1(n5674), .B2(n6775), .A(n103), .ZN(n3738) );
  OAI21_X2 U6929 ( .B1(n6779), .B2(n5674), .A(n38), .ZN(n3739) );
  OAI21_X2 U6930 ( .B1(n6660), .B2(net367593), .A(n1078), .ZN(n3740) );
  OAI21_X2 U6931 ( .B1(n6660), .B2(n6683), .A(n1045), .ZN(n3741) );
  OAI21_X2 U6932 ( .B1(n6660), .B2(n6686), .A(n1011), .ZN(n3742) );
  OAI21_X2 U6933 ( .B1(n6660), .B2(n6689), .A(n977), .ZN(n3743) );
  OAI21_X2 U6934 ( .B1(n6660), .B2(n6693), .A(n944), .ZN(n3744) );
  OAI21_X2 U6935 ( .B1(n6660), .B2(n6700), .A(n876), .ZN(n3746) );
  OAI21_X2 U6936 ( .B1(n6660), .B2(n6704), .A(n843), .ZN(n3747) );
  OAI21_X2 U6937 ( .B1(n6660), .B2(n6707), .A(n810), .ZN(n3748) );
  OAI21_X2 U6938 ( .B1(n6660), .B2(n6710), .A(n776), .ZN(n3749) );
  OAI21_X2 U6939 ( .B1(n6661), .B2(n6717), .A(n710), .ZN(n3750) );
  OAI21_X2 U6940 ( .B1(n6661), .B2(n6722), .A(n677), .ZN(n3751) );
  OAI21_X2 U6941 ( .B1(n6661), .B2(n6725), .A(n644), .ZN(n3752) );
  OAI21_X2 U6942 ( .B1(n6661), .B2(n6728), .A(n610), .ZN(n3753) );
  OAI21_X2 U6943 ( .B1(n6661), .B2(n6732), .A(n575), .ZN(n3754) );
  OAI21_X2 U6944 ( .B1(n6661), .B2(n6736), .A(n542), .ZN(n3755) );
  OAI21_X2 U6945 ( .B1(n6661), .B2(n6740), .A(n509), .ZN(n3756) );
  OAI21_X2 U6946 ( .B1(n6661), .B2(n6743), .A(n475), .ZN(n3757) );
  OAI21_X2 U6947 ( .B1(n6661), .B2(n439), .A(n441), .ZN(n3758) );
  OAI21_X2 U6948 ( .B1(n6661), .B2(n6749), .A(n408), .ZN(n3759) );
  OAI21_X2 U6949 ( .B1(n6661), .B2(n6752), .A(n342), .ZN(n3760) );
  AOI21_X2 U6950 ( .B1(drData[23]), .B2(n1158), .A(n13673), .ZN(n1183) );
  OAI21_X2 U6951 ( .B1(n6659), .B2(n6678), .A(n1110), .ZN(n3763) );
  OAI21_X2 U6952 ( .B1(n6659), .B2(n6713), .A(n742), .ZN(n3764) );
  OAI21_X2 U6953 ( .B1(n5675), .B2(net367215), .A(n374), .ZN(n3765) );
  OAI21_X2 U6954 ( .B1(n6659), .B2(n6758), .A(n273), .ZN(n3766) );
  OAI21_X2 U6955 ( .B1(n5675), .B2(n6761), .A(n238), .ZN(n3767) );
  OAI21_X2 U6956 ( .B1(n6659), .B2(n6765), .A(n205), .ZN(n3768) );
  OAI21_X2 U6957 ( .B1(n5675), .B2(n6768), .A(n171), .ZN(n3769) );
  OAI21_X2 U6958 ( .B1(n6659), .B2(n6775), .A(n102), .ZN(n3771) );
  OAI21_X2 U6959 ( .B1(n6659), .B2(net367593), .A(n1077), .ZN(n3773) );
  OAI21_X2 U6960 ( .B1(n6659), .B2(n6683), .A(n1044), .ZN(n3774) );
  OAI21_X2 U6961 ( .B1(n6659), .B2(n6686), .A(n1010), .ZN(n3775) );
  OAI21_X2 U6962 ( .B1(n6659), .B2(n6700), .A(n875), .ZN(n3779) );
  OAI21_X2 U6963 ( .B1(n6659), .B2(n6704), .A(n842), .ZN(n3780) );
  OAI21_X2 U6964 ( .B1(n6659), .B2(n6707), .A(n809), .ZN(n3781) );
  OAI21_X2 U6965 ( .B1(n6659), .B2(n6732), .A(n574), .ZN(n3787) );
  AOI21_X2 U6966 ( .B1(drData[22]), .B2(n1158), .A(n13673), .ZN(n1186) );
  OAI21_X2 U6967 ( .B1(n6658), .B2(n6678), .A(n1140), .ZN(n3796) );
  OAI21_X2 U6968 ( .B1(n6658), .B2(n6713), .A(n772), .ZN(n3797) );
  OAI21_X2 U6969 ( .B1(n6658), .B2(net367215), .A(n404), .ZN(n3798) );
  OAI21_X2 U6970 ( .B1(n5649), .B2(n6761), .A(n268), .ZN(n3800) );
  OAI21_X2 U6971 ( .B1(n6658), .B2(n6765), .A(n235), .ZN(n3801) );
  OAI21_X2 U6972 ( .B1(n5649), .B2(n6768), .A(n201), .ZN(n3802) );
  OAI21_X2 U6973 ( .B1(n6658), .B2(n6772), .A(n166), .ZN(n3803) );
  OAI21_X2 U6974 ( .B1(n6658), .B2(n6775), .A(n132), .ZN(n3804) );
  OAI21_X2 U6975 ( .B1(n6779), .B2(n5649), .A(n96), .ZN(n3805) );
  OAI21_X2 U6976 ( .B1(n6658), .B2(net367593), .A(n1107), .ZN(n3806) );
  OAI21_X2 U6977 ( .B1(n6658), .B2(n6686), .A(n1040), .ZN(n3808) );
  OAI21_X2 U6978 ( .B1(n6658), .B2(n6689), .A(n1006), .ZN(n3809) );
  OAI21_X2 U6979 ( .B1(n6658), .B2(n6700), .A(n905), .ZN(n3812) );
  OAI21_X2 U6980 ( .B1(n6658), .B2(n6704), .A(n872), .ZN(n3813) );
  OAI21_X2 U6981 ( .B1(n6658), .B2(n6707), .A(n839), .ZN(n3814) );
  OAI21_X2 U6982 ( .B1(n6658), .B2(n6717), .A(n739), .ZN(n3816) );
  OAI21_X2 U6983 ( .B1(n5649), .B2(n6732), .A(n604), .ZN(n3820) );
  AOI21_X2 U6984 ( .B1(drData[21]), .B2(n1158), .A(n13673), .ZN(n1189) );
  OAI21_X2 U6985 ( .B1(n6656), .B2(n6678), .A(n1139), .ZN(n3829) );
  OAI21_X2 U6986 ( .B1(n6656), .B2(n6713), .A(n771), .ZN(n3830) );
  OAI21_X2 U6987 ( .B1(n6657), .B2(net367215), .A(n403), .ZN(n3831) );
  OAI21_X2 U6988 ( .B1(n6657), .B2(n6758), .A(n302), .ZN(n3832) );
  OAI21_X2 U6989 ( .B1(n5650), .B2(n6761), .A(n267), .ZN(n3833) );
  OAI21_X2 U6990 ( .B1(n6656), .B2(n6765), .A(n234), .ZN(n3834) );
  OAI21_X2 U6991 ( .B1(n5650), .B2(n6768), .A(n200), .ZN(n3835) );
  OAI21_X2 U6992 ( .B1(n5650), .B2(n6772), .A(n165), .ZN(n3836) );
  OAI21_X2 U6993 ( .B1(n5650), .B2(n6775), .A(n131), .ZN(n3837) );
  OAI21_X2 U6994 ( .B1(n6779), .B2(n5650), .A(n94), .ZN(n3838) );
  OAI21_X2 U6995 ( .B1(n6656), .B2(net367593), .A(n1106), .ZN(n3839) );
  OAI21_X2 U6996 ( .B1(n6656), .B2(n6683), .A(n1073), .ZN(n3840) );
  OAI21_X2 U6997 ( .B1(n6656), .B2(n6686), .A(n1039), .ZN(n3841) );
  OAI21_X2 U6998 ( .B1(n6656), .B2(n6689), .A(n1005), .ZN(n3842) );
  OAI21_X2 U6999 ( .B1(n6656), .B2(n6693), .A(n972), .ZN(n3843) );
  OAI21_X2 U7000 ( .B1(n6656), .B2(n6697), .A(n938), .ZN(n3844) );
  OAI21_X2 U7001 ( .B1(n6656), .B2(n6700), .A(n904), .ZN(n3845) );
  OAI21_X2 U7002 ( .B1(n6656), .B2(n6704), .A(n871), .ZN(n3846) );
  OAI21_X2 U7003 ( .B1(n6656), .B2(n6707), .A(n838), .ZN(n3847) );
  OAI21_X2 U7004 ( .B1(n6656), .B2(n6710), .A(n804), .ZN(n3848) );
  OAI21_X2 U7005 ( .B1(n6657), .B2(n6717), .A(n738), .ZN(n3849) );
  OAI21_X2 U7006 ( .B1(n6657), .B2(n6722), .A(n705), .ZN(n3850) );
  OAI21_X2 U7007 ( .B1(n6657), .B2(n6725), .A(n672), .ZN(n3851) );
  OAI21_X2 U7008 ( .B1(n6657), .B2(n6728), .A(n638), .ZN(n3852) );
  OAI21_X2 U7009 ( .B1(n6657), .B2(n6732), .A(n603), .ZN(n3853) );
  OAI21_X2 U7010 ( .B1(n6657), .B2(n6736), .A(n570), .ZN(n3854) );
  OAI21_X2 U7011 ( .B1(n6657), .B2(n6740), .A(n537), .ZN(n3855) );
  OAI21_X2 U7012 ( .B1(n6657), .B2(n6743), .A(n503), .ZN(n3856) );
  OAI21_X2 U7013 ( .B1(n6657), .B2(n439), .A(n469), .ZN(n3857) );
  OAI21_X2 U7014 ( .B1(n6657), .B2(n6749), .A(n436), .ZN(n3858) );
  OAI21_X2 U7015 ( .B1(n6657), .B2(n6752), .A(n370), .ZN(n3859) );
  OAI21_X2 U7016 ( .B1(n6656), .B2(n6755), .A(n336), .ZN(n3860) );
  AOI21_X2 U7017 ( .B1(drData[20]), .B2(n1158), .A(n13673), .ZN(n1192) );
  OAI21_X2 U7018 ( .B1(n6655), .B2(n6678), .A(n1138), .ZN(n3862) );
  OAI21_X2 U7019 ( .B1(n6655), .B2(net367215), .A(n402), .ZN(n3864) );
  OAI21_X2 U7020 ( .B1(n5651), .B2(n6761), .A(n266), .ZN(n3866) );
  OAI21_X2 U7021 ( .B1(n6655), .B2(n6765), .A(n233), .ZN(n3867) );
  OAI21_X2 U7022 ( .B1(n6655), .B2(n6768), .A(n199), .ZN(n3868) );
  OAI21_X2 U7023 ( .B1(n6655), .B2(n6772), .A(n164), .ZN(n3869) );
  OAI21_X2 U7024 ( .B1(n5651), .B2(n6775), .A(n130), .ZN(n3870) );
  OAI21_X2 U7025 ( .B1(n6779), .B2(n5651), .A(n92), .ZN(n3871) );
  OAI21_X2 U7026 ( .B1(n5651), .B2(net367593), .A(n1105), .ZN(n3872) );
  OAI21_X2 U7027 ( .B1(n6655), .B2(n6683), .A(n1072), .ZN(n3873) );
  OAI21_X2 U7028 ( .B1(n6655), .B2(n6686), .A(n1038), .ZN(n3874) );
  OAI21_X2 U7029 ( .B1(n6655), .B2(n6689), .A(n1004), .ZN(n3875) );
  OAI21_X2 U7030 ( .B1(n6655), .B2(n6700), .A(n903), .ZN(n3878) );
  OAI21_X2 U7031 ( .B1(n6655), .B2(n6704), .A(n870), .ZN(n3879) );
  OAI21_X2 U7032 ( .B1(n6655), .B2(n6707), .A(n837), .ZN(n3880) );
  OAI21_X2 U7033 ( .B1(n5651), .B2(n6710), .A(n803), .ZN(n3881) );
  OAI21_X2 U7034 ( .B1(n6655), .B2(n6717), .A(n737), .ZN(n3882) );
  OAI21_X2 U7035 ( .B1(n6655), .B2(n6722), .A(n704), .ZN(n3883) );
  OAI21_X2 U7036 ( .B1(n6655), .B2(n6725), .A(n671), .ZN(n3884) );
  OAI21_X2 U7037 ( .B1(n6655), .B2(n6728), .A(n637), .ZN(n3885) );
  OAI21_X2 U7038 ( .B1(n6655), .B2(n6732), .A(n602), .ZN(n3886) );
  OAI21_X2 U7039 ( .B1(n6655), .B2(n6736), .A(n569), .ZN(n3887) );
  OAI21_X2 U7040 ( .B1(n6655), .B2(n6740), .A(n536), .ZN(n3888) );
  OAI21_X2 U7041 ( .B1(n6655), .B2(n6743), .A(n502), .ZN(n3889) );
  OAI21_X2 U7042 ( .B1(n6655), .B2(n439), .A(n468), .ZN(n3890) );
  OAI21_X2 U7043 ( .B1(n6655), .B2(n6749), .A(n435), .ZN(n3891) );
  OAI21_X2 U7044 ( .B1(n6655), .B2(n6752), .A(n369), .ZN(n3892) );
  OAI21_X2 U7045 ( .B1(n5651), .B2(n6755), .A(n335), .ZN(n3893) );
  AOI21_X2 U7046 ( .B1(drData[19]), .B2(n1158), .A(n13673), .ZN(n1195) );
  OAI21_X2 U7047 ( .B1(n6653), .B2(n6679), .A(n1137), .ZN(n3895) );
  OAI21_X2 U7048 ( .B1(n6653), .B2(n6714), .A(n769), .ZN(n3896) );
  OAI21_X2 U7049 ( .B1(n6654), .B2(net367217), .A(n401), .ZN(n3897) );
  OAI21_X2 U7050 ( .B1(n6653), .B2(n6759), .A(n300), .ZN(n3898) );
  OAI21_X2 U7051 ( .B1(n5652), .B2(n6762), .A(n265), .ZN(n3899) );
  OAI21_X2 U7052 ( .B1(n6653), .B2(n6766), .A(n232), .ZN(n3900) );
  OAI21_X2 U7053 ( .B1(n5652), .B2(n6769), .A(n198), .ZN(n3901) );
  OAI21_X2 U7054 ( .B1(n6654), .B2(n6773), .A(n163), .ZN(n3902) );
  OAI21_X2 U7055 ( .B1(n5652), .B2(n6776), .A(n129), .ZN(n3903) );
  OAI21_X2 U7056 ( .B1(n6780), .B2(n5652), .A(n90), .ZN(n3904) );
  OAI21_X2 U7057 ( .B1(n6653), .B2(net367595), .A(n1104), .ZN(n3905) );
  OAI21_X2 U7058 ( .B1(n6653), .B2(n6684), .A(n1071), .ZN(n3906) );
  OAI21_X2 U7059 ( .B1(n6653), .B2(n6687), .A(n1037), .ZN(n3907) );
  OAI21_X2 U7060 ( .B1(n6653), .B2(n6690), .A(n1003), .ZN(n3908) );
  OAI21_X2 U7061 ( .B1(n6653), .B2(n6694), .A(n970), .ZN(n3909) );
  OAI21_X2 U7062 ( .B1(n6653), .B2(n6698), .A(n936), .ZN(n3910) );
  OAI21_X2 U7063 ( .B1(n6653), .B2(n6701), .A(n902), .ZN(n3911) );
  OAI21_X2 U7064 ( .B1(n6653), .B2(n6705), .A(n869), .ZN(n3912) );
  OAI21_X2 U7065 ( .B1(n6653), .B2(n6708), .A(n836), .ZN(n3913) );
  OAI21_X2 U7066 ( .B1(n6653), .B2(n6711), .A(n802), .ZN(n3914) );
  OAI21_X2 U7067 ( .B1(n6654), .B2(n6718), .A(n736), .ZN(n3915) );
  OAI21_X2 U7068 ( .B1(n6654), .B2(n6723), .A(n703), .ZN(n3916) );
  OAI21_X2 U7069 ( .B1(n6654), .B2(n6726), .A(n670), .ZN(n3917) );
  OAI21_X2 U7070 ( .B1(n6654), .B2(n6729), .A(n636), .ZN(n3918) );
  OAI21_X2 U7071 ( .B1(n6654), .B2(n6733), .A(n601), .ZN(n3919) );
  OAI21_X2 U7072 ( .B1(n6654), .B2(n6737), .A(n568), .ZN(n3920) );
  OAI21_X2 U7073 ( .B1(n6654), .B2(n6741), .A(n535), .ZN(n3921) );
  OAI21_X2 U7074 ( .B1(n6654), .B2(n6744), .A(n501), .ZN(n3922) );
  OAI21_X2 U7075 ( .B1(n6654), .B2(n6750), .A(n434), .ZN(n3924) );
  AOI21_X2 U7076 ( .B1(drData[18]), .B2(n1158), .A(n13673), .ZN(n1198) );
  OAI21_X2 U7077 ( .B1(n6651), .B2(n6679), .A(n1136), .ZN(n3928) );
  OAI21_X2 U7078 ( .B1(n6651), .B2(n6714), .A(n768), .ZN(n3929) );
  OAI21_X2 U7079 ( .B1(n5653), .B2(n6759), .A(n299), .ZN(n3931) );
  OAI21_X2 U7080 ( .B1(n6651), .B2(n6762), .A(n264), .ZN(n3932) );
  OAI21_X2 U7081 ( .B1(n6651), .B2(n6766), .A(n231), .ZN(n3933) );
  OAI21_X2 U7082 ( .B1(n5653), .B2(n6769), .A(n197), .ZN(n3934) );
  OAI21_X2 U7083 ( .B1(n6652), .B2(n6773), .A(n162), .ZN(n3935) );
  OAI21_X2 U7084 ( .B1(n5653), .B2(n6776), .A(n128), .ZN(n3936) );
  OAI21_X2 U7085 ( .B1(n6780), .B2(n5653), .A(n88), .ZN(n3937) );
  OAI21_X2 U7086 ( .B1(n6651), .B2(n6684), .A(n1070), .ZN(n3939) );
  OAI21_X2 U7087 ( .B1(n6651), .B2(n6687), .A(n1036), .ZN(n3940) );
  OAI21_X2 U7088 ( .B1(n6651), .B2(n6690), .A(n1002), .ZN(n3941) );
  OAI21_X2 U7089 ( .B1(n6651), .B2(n6694), .A(n969), .ZN(n3942) );
  OAI21_X2 U7090 ( .B1(n6651), .B2(n6698), .A(n935), .ZN(n3943) );
  OAI21_X2 U7091 ( .B1(n6651), .B2(n6701), .A(n901), .ZN(n3944) );
  OAI21_X2 U7092 ( .B1(n6651), .B2(n6705), .A(n868), .ZN(n3945) );
  OAI21_X2 U7093 ( .B1(n6651), .B2(n6711), .A(n801), .ZN(n3947) );
  OAI21_X2 U7094 ( .B1(n6652), .B2(n6718), .A(n735), .ZN(n3948) );
  OAI21_X2 U7095 ( .B1(n6652), .B2(n6723), .A(n702), .ZN(n3949) );
  OAI21_X2 U7096 ( .B1(n6652), .B2(n6726), .A(n669), .ZN(n3950) );
  OAI21_X2 U7097 ( .B1(n6652), .B2(n6729), .A(n635), .ZN(n3951) );
  OAI21_X2 U7098 ( .B1(n6652), .B2(n6733), .A(n600), .ZN(n3952) );
  OAI21_X2 U7099 ( .B1(n6652), .B2(n6737), .A(n567), .ZN(n3953) );
  OAI21_X2 U7100 ( .B1(n6652), .B2(n6744), .A(n500), .ZN(n3955) );
  OAI21_X2 U7101 ( .B1(n6652), .B2(n6747), .A(n466), .ZN(n3956) );
  OAI21_X2 U7102 ( .B1(n6652), .B2(n6750), .A(n433), .ZN(n3957) );
  OAI21_X2 U7103 ( .B1(n6652), .B2(n6753), .A(n367), .ZN(n3958) );
  OAI21_X2 U7104 ( .B1(n5653), .B2(n6756), .A(n333), .ZN(n3959) );
  AOI21_X2 U7105 ( .B1(drData[17]), .B2(n1158), .A(n13673), .ZN(n1201) );
  OAI21_X2 U7106 ( .B1(n6649), .B2(n6714), .A(n767), .ZN(n3962) );
  OAI21_X2 U7107 ( .B1(n5654), .B2(n6759), .A(n298), .ZN(n3964) );
  OAI21_X2 U7108 ( .B1(n5654), .B2(n6762), .A(n263), .ZN(n3965) );
  OAI21_X2 U7109 ( .B1(n6650), .B2(n6766), .A(n230), .ZN(n3966) );
  OAI21_X2 U7110 ( .B1(n5654), .B2(n6769), .A(n196), .ZN(n3967) );
  OAI21_X2 U7111 ( .B1(n6649), .B2(n6773), .A(n161), .ZN(n3968) );
  OAI21_X2 U7112 ( .B1(n5654), .B2(n6776), .A(n127), .ZN(n3969) );
  OAI21_X2 U7113 ( .B1(n6780), .B2(n5654), .A(n86), .ZN(n3970) );
  OAI21_X2 U7114 ( .B1(n6649), .B2(net367595), .A(n1102), .ZN(n3971) );
  OAI21_X2 U7115 ( .B1(n6649), .B2(n6684), .A(n1069), .ZN(n3972) );
  OAI21_X2 U7116 ( .B1(n6649), .B2(n6687), .A(n1035), .ZN(n3973) );
  OAI21_X2 U7117 ( .B1(n6649), .B2(n6690), .A(n1001), .ZN(n3974) );
  OAI21_X2 U7118 ( .B1(n6649), .B2(n6694), .A(n968), .ZN(n3975) );
  OAI21_X2 U7119 ( .B1(n6649), .B2(n6698), .A(n934), .ZN(n3976) );
  OAI21_X2 U7120 ( .B1(n6649), .B2(n6705), .A(n867), .ZN(n3978) );
  OAI21_X2 U7121 ( .B1(n6649), .B2(n6711), .A(n800), .ZN(n3980) );
  OAI21_X2 U7122 ( .B1(n6650), .B2(n6718), .A(n734), .ZN(n3981) );
  OAI21_X2 U7123 ( .B1(n6650), .B2(n6723), .A(n701), .ZN(n3982) );
  OAI21_X2 U7124 ( .B1(n6650), .B2(n6726), .A(n668), .ZN(n3983) );
  OAI21_X2 U7125 ( .B1(n6650), .B2(n6729), .A(n634), .ZN(n3984) );
  OAI21_X2 U7126 ( .B1(n6650), .B2(n6737), .A(n566), .ZN(n3986) );
  OAI21_X2 U7127 ( .B1(n6650), .B2(n6744), .A(n499), .ZN(n3988) );
  OAI21_X2 U7128 ( .B1(n6650), .B2(n6747), .A(n465), .ZN(n3989) );
  OAI21_X2 U7129 ( .B1(n6650), .B2(n6750), .A(n432), .ZN(n3990) );
  OAI21_X2 U7130 ( .B1(n6650), .B2(n6753), .A(n366), .ZN(n3991) );
  OAI21_X2 U7131 ( .B1(n6649), .B2(n6756), .A(n332), .ZN(n3992) );
  AOI21_X2 U7132 ( .B1(drData[16]), .B2(n1158), .A(n13673), .ZN(n1204) );
  OAI21_X2 U7133 ( .B1(n6647), .B2(n1109), .A(n1134), .ZN(n3994) );
  OAI21_X2 U7134 ( .B1(n6647), .B2(n741), .A(n766), .ZN(n3995) );
  OAI21_X2 U7135 ( .B1(n6648), .B2(net367215), .A(n398), .ZN(n3996) );
  OAI21_X2 U7136 ( .B1(n6648), .B2(n6760), .A(n297), .ZN(n3997) );
  OAI21_X2 U7137 ( .B1(n5655), .B2(n237), .A(n262), .ZN(n3998) );
  OAI21_X2 U7138 ( .B1(n6647), .B2(n6767), .A(n229), .ZN(n3999) );
  OAI21_X2 U7139 ( .B1(n5655), .B2(n6770), .A(n195), .ZN(n4000) );
  OAI21_X2 U7140 ( .B1(n6648), .B2(n6774), .A(n160), .ZN(n4001) );
  OAI21_X2 U7141 ( .B1(n5655), .B2(n6777), .A(n126), .ZN(n4002) );
  OAI21_X2 U7142 ( .B1(n34), .B2(n5655), .A(n84), .ZN(n4003) );
  OAI21_X2 U7143 ( .B1(n6647), .B2(net367597), .A(n1101), .ZN(n4004) );
  OAI21_X2 U7144 ( .B1(n6647), .B2(n1043), .A(n1068), .ZN(n4005) );
  OAI21_X2 U7145 ( .B1(n6647), .B2(n6688), .A(n1034), .ZN(n4006) );
  OAI21_X2 U7146 ( .B1(n6647), .B2(n6691), .A(n1000), .ZN(n4007) );
  OAI21_X2 U7147 ( .B1(n6647), .B2(n6702), .A(n899), .ZN(n4010) );
  OAI21_X2 U7148 ( .B1(n6647), .B2(n6706), .A(n866), .ZN(n4011) );
  OAI21_X2 U7149 ( .B1(n6647), .B2(n6709), .A(n833), .ZN(n4012) );
  OAI21_X2 U7150 ( .B1(n6647), .B2(n6712), .A(n799), .ZN(n4013) );
  OAI21_X2 U7151 ( .B1(n6648), .B2(n708), .A(n733), .ZN(n4014) );
  OAI21_X2 U7152 ( .B1(n6648), .B2(n6723), .A(n700), .ZN(n4015) );
  OAI21_X2 U7153 ( .B1(n6648), .B2(n6727), .A(n667), .ZN(n4016) );
  OAI21_X2 U7154 ( .B1(n6648), .B2(n6730), .A(n633), .ZN(n4017) );
  OAI21_X2 U7155 ( .B1(n6648), .B2(n6734), .A(n598), .ZN(n4018) );
  OAI21_X2 U7156 ( .B1(n6648), .B2(n540), .A(n565), .ZN(n4019) );
  OAI21_X2 U7157 ( .B1(n6648), .B2(n507), .A(n532), .ZN(n4020) );
  OAI21_X2 U7158 ( .B1(n6648), .B2(n6745), .A(n498), .ZN(n4021) );
  OAI21_X2 U7159 ( .B1(n6648), .B2(n6747), .A(n464), .ZN(n4022) );
  OAI21_X2 U7160 ( .B1(n6648), .B2(n6751), .A(n431), .ZN(n4023) );
  OAI21_X2 U7161 ( .B1(n6648), .B2(n6752), .A(n365), .ZN(n4024) );
  OAI21_X2 U7162 ( .B1(n6645), .B2(n1109), .A(n1133), .ZN(n4027) );
  OAI21_X2 U7163 ( .B1(n6645), .B2(n741), .A(n765), .ZN(n4028) );
  OAI21_X2 U7164 ( .B1(n6646), .B2(n373), .A(n397), .ZN(n4029) );
  OAI21_X2 U7165 ( .B1(n6645), .B2(n6760), .A(n296), .ZN(n4030) );
  OAI21_X2 U7166 ( .B1(n5656), .B2(n6762), .A(n261), .ZN(n4031) );
  OAI21_X2 U7167 ( .B1(n6646), .B2(n6767), .A(n228), .ZN(n4032) );
  OAI21_X2 U7168 ( .B1(n5656), .B2(n6770), .A(n194), .ZN(n4033) );
  OAI21_X2 U7169 ( .B1(n6645), .B2(n6774), .A(n159), .ZN(n4034) );
  OAI21_X2 U7170 ( .B1(n5656), .B2(n6777), .A(n125), .ZN(n4035) );
  OAI21_X2 U7171 ( .B1(n34), .B2(n5656), .A(n82), .ZN(n4036) );
  OAI21_X2 U7172 ( .B1(n6645), .B2(net367597), .A(n1100), .ZN(n4037) );
  OAI21_X2 U7173 ( .B1(n6645), .B2(n1043), .A(n1067), .ZN(n4038) );
  OAI21_X2 U7174 ( .B1(n6645), .B2(n6688), .A(n1033), .ZN(n4039) );
  OAI21_X2 U7175 ( .B1(n6645), .B2(n6691), .A(n999), .ZN(n4040) );
  OAI21_X2 U7176 ( .B1(n6645), .B2(n942), .A(n966), .ZN(n4041) );
  OAI21_X2 U7177 ( .B1(n6645), .B2(n6699), .A(n932), .ZN(n4042) );
  OAI21_X2 U7178 ( .B1(n6645), .B2(n6702), .A(n898), .ZN(n4043) );
  OAI21_X2 U7179 ( .B1(n6645), .B2(n6706), .A(n865), .ZN(n4044) );
  OAI21_X2 U7180 ( .B1(n6645), .B2(n6709), .A(n832), .ZN(n4045) );
  OAI21_X2 U7181 ( .B1(n6645), .B2(n6712), .A(n798), .ZN(n4046) );
  OAI21_X2 U7182 ( .B1(n6646), .B2(n708), .A(n732), .ZN(n4047) );
  OAI21_X2 U7183 ( .B1(n6646), .B2(n675), .A(n699), .ZN(n4048) );
  OAI21_X2 U7184 ( .B1(n6646), .B2(n6727), .A(n666), .ZN(n4049) );
  OAI21_X2 U7185 ( .B1(n6646), .B2(n6730), .A(n632), .ZN(n4050) );
  OAI21_X2 U7186 ( .B1(n6646), .B2(n6734), .A(n597), .ZN(n4051) );
  OAI21_X2 U7187 ( .B1(n6646), .B2(n540), .A(n564), .ZN(n4052) );
  OAI21_X2 U7188 ( .B1(n6646), .B2(n507), .A(n531), .ZN(n4053) );
  OAI21_X2 U7189 ( .B1(n6646), .B2(n6745), .A(n497), .ZN(n4054) );
  OAI21_X2 U7190 ( .B1(n6646), .B2(n6748), .A(n463), .ZN(n4055) );
  OAI21_X2 U7191 ( .B1(n6646), .B2(n6751), .A(n430), .ZN(n4056) );
  OAI21_X2 U7192 ( .B1(n6646), .B2(n6753), .A(n364), .ZN(n4057) );
  OAI21_X2 U7193 ( .B1(n5656), .B2(n6757), .A(n330), .ZN(n4058) );
  OAI21_X2 U7194 ( .B1(n6644), .B2(n6679), .A(n1132), .ZN(n4060) );
  OAI21_X2 U7195 ( .B1(n6644), .B2(n6714), .A(n764), .ZN(n4061) );
  OAI21_X2 U7196 ( .B1(n5657), .B2(net367221), .A(n396), .ZN(n4062) );
  OAI21_X2 U7197 ( .B1(n6644), .B2(n6760), .A(n295), .ZN(n4063) );
  OAI21_X2 U7198 ( .B1(n5657), .B2(n6761), .A(n260), .ZN(n4064) );
  OAI21_X2 U7199 ( .B1(n6644), .B2(n6767), .A(n227), .ZN(n4065) );
  OAI21_X2 U7200 ( .B1(n5657), .B2(n6770), .A(n193), .ZN(n4066) );
  OAI21_X2 U7201 ( .B1(n6644), .B2(n6774), .A(n158), .ZN(n4067) );
  OAI21_X2 U7202 ( .B1(n5657), .B2(n6777), .A(n124), .ZN(n4068) );
  OAI21_X2 U7203 ( .B1(n6779), .B2(n5657), .A(n80), .ZN(n4069) );
  OAI21_X2 U7204 ( .B1(n6644), .B2(net367597), .A(n1099), .ZN(n4070) );
  OAI21_X2 U7205 ( .B1(n6644), .B2(n6685), .A(n1066), .ZN(n4071) );
  OAI21_X2 U7206 ( .B1(n6644), .B2(n6688), .A(n1032), .ZN(n4072) );
  OAI21_X2 U7207 ( .B1(n6644), .B2(n6691), .A(n998), .ZN(n4073) );
  OAI21_X2 U7208 ( .B1(n6644), .B2(n6693), .A(n965), .ZN(n4074) );
  OAI21_X2 U7209 ( .B1(n6644), .B2(n6699), .A(n931), .ZN(n4075) );
  OAI21_X2 U7210 ( .B1(n6644), .B2(n6702), .A(n897), .ZN(n4076) );
  OAI21_X2 U7211 ( .B1(n6644), .B2(n6706), .A(n864), .ZN(n4077) );
  OAI21_X2 U7212 ( .B1(n6644), .B2(n6709), .A(n831), .ZN(n4078) );
  OAI21_X2 U7213 ( .B1(n6644), .B2(n6712), .A(n797), .ZN(n4079) );
  OAI21_X2 U7214 ( .B1(n5657), .B2(n6719), .A(n731), .ZN(n4080) );
  OAI21_X2 U7215 ( .B1(n6644), .B2(n6724), .A(n698), .ZN(n4081) );
  OAI21_X2 U7216 ( .B1(n6644), .B2(n6727), .A(n665), .ZN(n4082) );
  OAI21_X2 U7217 ( .B1(n6644), .B2(n6730), .A(n631), .ZN(n4083) );
  OAI21_X2 U7218 ( .B1(n5657), .B2(n6738), .A(n563), .ZN(n4085) );
  OAI21_X2 U7219 ( .B1(n6644), .B2(n6742), .A(n530), .ZN(n4086) );
  OAI21_X2 U7220 ( .B1(n6644), .B2(n6745), .A(n496), .ZN(n4087) );
  OAI21_X2 U7221 ( .B1(n6644), .B2(n6748), .A(n462), .ZN(n4088) );
  OAI21_X2 U7222 ( .B1(n6644), .B2(n6751), .A(n429), .ZN(n4089) );
  OAI21_X2 U7223 ( .B1(n6644), .B2(n340), .A(n363), .ZN(n4090) );
  OAI21_X2 U7224 ( .B1(n5657), .B2(n6757), .A(n329), .ZN(n4091) );
  OAI21_X2 U7225 ( .B1(n6642), .B2(n1109), .A(n1131), .ZN(n4093) );
  OAI21_X2 U7226 ( .B1(n6642), .B2(n741), .A(n763), .ZN(n4094) );
  OAI21_X2 U7227 ( .B1(n6643), .B2(n373), .A(n395), .ZN(n4095) );
  OAI21_X2 U7228 ( .B1(n6642), .B2(n6760), .A(n294), .ZN(n4096) );
  OAI21_X2 U7229 ( .B1(n5658), .B2(n237), .A(n259), .ZN(n4097) );
  OAI21_X2 U7230 ( .B1(n6643), .B2(n6767), .A(n226), .ZN(n4098) );
  OAI21_X2 U7231 ( .B1(n5658), .B2(n6770), .A(n192), .ZN(n4099) );
  OAI21_X2 U7232 ( .B1(n6642), .B2(n6774), .A(n157), .ZN(n4100) );
  OAI21_X2 U7233 ( .B1(n5658), .B2(n6777), .A(n123), .ZN(n4101) );
  OAI21_X2 U7234 ( .B1(n34), .B2(n5658), .A(n78), .ZN(n4102) );
  OAI21_X2 U7235 ( .B1(n6642), .B2(net367597), .A(n1098), .ZN(n4103) );
  OAI21_X2 U7236 ( .B1(n6642), .B2(n1043), .A(n1065), .ZN(n4104) );
  OAI21_X2 U7237 ( .B1(n6642), .B2(n6688), .A(n1031), .ZN(n4105) );
  OAI21_X2 U7238 ( .B1(n6642), .B2(n6691), .A(n997), .ZN(n4106) );
  OAI21_X2 U7239 ( .B1(n6642), .B2(n942), .A(n964), .ZN(n4107) );
  OAI21_X2 U7240 ( .B1(n6642), .B2(n6699), .A(n930), .ZN(n4108) );
  OAI21_X2 U7241 ( .B1(n6642), .B2(n6702), .A(n896), .ZN(n4109) );
  OAI21_X2 U7242 ( .B1(n6642), .B2(n6706), .A(n863), .ZN(n4110) );
  OAI21_X2 U7243 ( .B1(n6642), .B2(n6709), .A(n830), .ZN(n4111) );
  OAI21_X2 U7244 ( .B1(n6642), .B2(n6712), .A(n796), .ZN(n4112) );
  OAI21_X2 U7245 ( .B1(n6643), .B2(n708), .A(n730), .ZN(n4113) );
  OAI21_X2 U7246 ( .B1(n6643), .B2(n675), .A(n697), .ZN(n4114) );
  OAI21_X2 U7247 ( .B1(n6643), .B2(n6727), .A(n664), .ZN(n4115) );
  OAI21_X2 U7248 ( .B1(n6643), .B2(n6730), .A(n630), .ZN(n4116) );
  OAI21_X2 U7249 ( .B1(n6643), .B2(n6734), .A(n595), .ZN(n4117) );
  OAI21_X2 U7250 ( .B1(n6643), .B2(n540), .A(n562), .ZN(n4118) );
  OAI21_X2 U7251 ( .B1(n6643), .B2(n507), .A(n529), .ZN(n4119) );
  OAI21_X2 U7252 ( .B1(n6643), .B2(n6745), .A(n495), .ZN(n4120) );
  OAI21_X2 U7253 ( .B1(n6643), .B2(n439), .A(n461), .ZN(n4121) );
  OAI21_X2 U7254 ( .B1(n6643), .B2(n6751), .A(n428), .ZN(n4122) );
  OAI21_X2 U7255 ( .B1(n6643), .B2(n6753), .A(n362), .ZN(n4123) );
  OAI21_X2 U7256 ( .B1(n5658), .B2(n6757), .A(n328), .ZN(n4124) );
  OAI21_X2 U7257 ( .B1(n6640), .B2(n6680), .A(n1129), .ZN(n4126) );
  OAI21_X2 U7258 ( .B1(n6640), .B2(n6715), .A(n761), .ZN(n4127) );
  OAI21_X2 U7259 ( .B1(n6641), .B2(n373), .A(n393), .ZN(n4128) );
  OAI21_X2 U7260 ( .B1(n6640), .B2(n6760), .A(n292), .ZN(n4129) );
  OAI21_X2 U7261 ( .B1(n5660), .B2(n6763), .A(n257), .ZN(n4130) );
  OAI21_X2 U7262 ( .B1(n6641), .B2(n6767), .A(n224), .ZN(n4131) );
  OAI21_X2 U7263 ( .B1(n5660), .B2(n6770), .A(n190), .ZN(n4132) );
  OAI21_X2 U7264 ( .B1(n6640), .B2(n6774), .A(n155), .ZN(n4133) );
  OAI21_X2 U7265 ( .B1(n5660), .B2(n6777), .A(n121), .ZN(n4134) );
  OAI21_X2 U7266 ( .B1(n6781), .B2(n5660), .A(n74), .ZN(n4135) );
  OAI21_X2 U7267 ( .B1(n6640), .B2(net367597), .A(n1096), .ZN(n4136) );
  OAI21_X2 U7268 ( .B1(n6640), .B2(n6683), .A(n1063), .ZN(n4137) );
  OAI21_X2 U7269 ( .B1(n6640), .B2(n6688), .A(n1029), .ZN(n4138) );
  OAI21_X2 U7270 ( .B1(n6640), .B2(n6691), .A(n995), .ZN(n4139) );
  OAI21_X2 U7271 ( .B1(n6640), .B2(n942), .A(n962), .ZN(n4140) );
  OAI21_X2 U7272 ( .B1(n6640), .B2(n6699), .A(n928), .ZN(n4141) );
  OAI21_X2 U7273 ( .B1(n6640), .B2(n6702), .A(n894), .ZN(n4142) );
  OAI21_X2 U7274 ( .B1(n6640), .B2(n6706), .A(n861), .ZN(n4143) );
  OAI21_X2 U7275 ( .B1(n6640), .B2(n6709), .A(n828), .ZN(n4144) );
  OAI21_X2 U7276 ( .B1(n6640), .B2(n6712), .A(n794), .ZN(n4145) );
  OAI21_X2 U7277 ( .B1(n6641), .B2(n708), .A(n728), .ZN(n4146) );
  OAI21_X2 U7278 ( .B1(n6641), .B2(n675), .A(n695), .ZN(n4147) );
  OAI21_X2 U7279 ( .B1(n6641), .B2(n6727), .A(n662), .ZN(n4148) );
  OAI21_X2 U7280 ( .B1(n6641), .B2(n6730), .A(n628), .ZN(n4149) );
  OAI21_X2 U7281 ( .B1(n6641), .B2(n6734), .A(n593), .ZN(n4150) );
  OAI21_X2 U7282 ( .B1(n6641), .B2(n540), .A(n560), .ZN(n4151) );
  OAI21_X2 U7283 ( .B1(n6641), .B2(n507), .A(n527), .ZN(n4152) );
  OAI21_X2 U7284 ( .B1(n6641), .B2(n6745), .A(n493), .ZN(n4153) );
  OAI21_X2 U7285 ( .B1(n6641), .B2(n439), .A(n459), .ZN(n4154) );
  OAI21_X2 U7286 ( .B1(n6641), .B2(n6751), .A(n426), .ZN(n4155) );
  OAI21_X2 U7287 ( .B1(n6641), .B2(n6752), .A(n360), .ZN(n4156) );
  OAI21_X2 U7288 ( .B1(n5660), .B2(n6757), .A(n326), .ZN(n4157) );
  OAI21_X2 U7289 ( .B1(n6638), .B2(n6714), .A(n760), .ZN(n4160) );
  OAI21_X2 U7290 ( .B1(n6639), .B2(net367217), .A(n392), .ZN(n4161) );
  OAI21_X2 U7291 ( .B1(n5661), .B2(n6759), .A(n291), .ZN(n4162) );
  OAI21_X2 U7292 ( .B1(n5661), .B2(n6762), .A(n256), .ZN(n4163) );
  OAI21_X2 U7293 ( .B1(n6639), .B2(n6766), .A(n223), .ZN(n4164) );
  OAI21_X2 U7294 ( .B1(n5661), .B2(n6769), .A(n189), .ZN(n4165) );
  OAI21_X2 U7295 ( .B1(n6638), .B2(n6773), .A(n154), .ZN(n4166) );
  OAI21_X2 U7296 ( .B1(n6780), .B2(n5661), .A(n72), .ZN(n4168) );
  OAI21_X2 U7297 ( .B1(n6638), .B2(net367595), .A(n1095), .ZN(n4169) );
  OAI21_X2 U7298 ( .B1(n6638), .B2(n6684), .A(n1062), .ZN(n4170) );
  OAI21_X2 U7299 ( .B1(n6638), .B2(n6687), .A(n1028), .ZN(n4171) );
  OAI21_X2 U7300 ( .B1(n6638), .B2(n6690), .A(n994), .ZN(n4172) );
  OAI21_X2 U7301 ( .B1(n6638), .B2(n6694), .A(n961), .ZN(n4173) );
  OAI21_X2 U7302 ( .B1(n6638), .B2(n6698), .A(n927), .ZN(n4174) );
  OAI21_X2 U7303 ( .B1(n6639), .B2(n6718), .A(n727), .ZN(n4179) );
  OAI21_X2 U7304 ( .B1(n6639), .B2(n6723), .A(n694), .ZN(n4180) );
  INV_X4 U7305 ( .A(n6955), .ZN(n6920) );
  OAI21_X2 U7306 ( .B1(n6639), .B2(n6726), .A(n661), .ZN(n4181) );
  OAI21_X2 U7307 ( .B1(n6639), .B2(n6729), .A(n627), .ZN(n4182) );
  OAI21_X2 U7308 ( .B1(n6639), .B2(n6737), .A(n559), .ZN(n4184) );
  OAI21_X2 U7309 ( .B1(n6639), .B2(n6744), .A(n492), .ZN(n4186) );
  OAI21_X2 U7310 ( .B1(n6639), .B2(n6747), .A(n458), .ZN(n4187) );
  OAI21_X2 U7311 ( .B1(n6639), .B2(n6750), .A(n425), .ZN(n4188) );
  INV_X4 U7312 ( .A(n6956), .ZN(n6932) );
  OAI21_X2 U7313 ( .B1(n6639), .B2(n6753), .A(n359), .ZN(n4189) );
  OAI21_X2 U7314 ( .B1(n6638), .B2(n6756), .A(n325), .ZN(n4190) );
  OAI21_X2 U7315 ( .B1(n6636), .B2(n1109), .A(n1127), .ZN(n4192) );
  OAI21_X2 U7316 ( .B1(n6636), .B2(n741), .A(n759), .ZN(n4193) );
  OAI21_X2 U7317 ( .B1(n6637), .B2(net367217), .A(n391), .ZN(n4194) );
  OAI21_X2 U7318 ( .B1(n6637), .B2(n6760), .A(n290), .ZN(n4195) );
  OAI21_X2 U7319 ( .B1(n5662), .B2(n237), .A(n255), .ZN(n4196) );
  OAI21_X2 U7320 ( .B1(n6636), .B2(n6767), .A(n222), .ZN(n4197) );
  OAI21_X2 U7321 ( .B1(n5662), .B2(n6770), .A(n188), .ZN(n4198) );
  OAI21_X2 U7322 ( .B1(n6637), .B2(n6774), .A(n153), .ZN(n4199) );
  OAI21_X2 U7323 ( .B1(n5662), .B2(n6777), .A(n119), .ZN(n4200) );
  OAI21_X2 U7324 ( .B1(n34), .B2(n5662), .A(n70), .ZN(n4201) );
  OAI21_X2 U7325 ( .B1(n6636), .B2(net367597), .A(n1094), .ZN(n4202) );
  OAI21_X2 U7326 ( .B1(n6636), .B2(n1043), .A(n1061), .ZN(n4203) );
  OAI21_X2 U7327 ( .B1(n6636), .B2(n6688), .A(n1027), .ZN(n4204) );
  OAI21_X2 U7328 ( .B1(n6636), .B2(n6691), .A(n993), .ZN(n4205) );
  OAI21_X2 U7329 ( .B1(n6636), .B2(n942), .A(n960), .ZN(n4206) );
  OAI21_X2 U7330 ( .B1(n6636), .B2(n6702), .A(n892), .ZN(n4208) );
  OAI21_X2 U7331 ( .B1(n6636), .B2(n6706), .A(n859), .ZN(n4209) );
  OAI21_X2 U7332 ( .B1(n6636), .B2(n6709), .A(n826), .ZN(n4210) );
  OAI21_X2 U7333 ( .B1(n6636), .B2(n6712), .A(n792), .ZN(n4211) );
  OAI21_X2 U7334 ( .B1(n6637), .B2(n708), .A(n726), .ZN(n4212) );
  OAI21_X2 U7335 ( .B1(n6637), .B2(n6722), .A(n693), .ZN(n4213) );
  OAI21_X2 U7336 ( .B1(n6637), .B2(n6727), .A(n660), .ZN(n4214) );
  OAI21_X2 U7337 ( .B1(n6637), .B2(n6730), .A(n626), .ZN(n4215) );
  OAI21_X2 U7338 ( .B1(n6637), .B2(n6734), .A(n591), .ZN(n4216) );
  OAI21_X2 U7339 ( .B1(n6637), .B2(n540), .A(n558), .ZN(n4217) );
  OAI21_X2 U7340 ( .B1(n6637), .B2(n507), .A(n525), .ZN(n4218) );
  OAI21_X2 U7341 ( .B1(n6637), .B2(n6745), .A(n491), .ZN(n4219) );
  OAI21_X2 U7342 ( .B1(n6637), .B2(n6748), .A(n457), .ZN(n4220) );
  OAI21_X2 U7343 ( .B1(n6637), .B2(n6751), .A(n424), .ZN(n4221) );
  OAI21_X2 U7344 ( .B1(n6637), .B2(n6752), .A(n358), .ZN(n4222) );
  OAI21_X2 U7345 ( .B1(n5662), .B2(n6757), .A(n324), .ZN(n4223) );
  OAI21_X2 U7346 ( .B1(n6634), .B2(n1109), .A(n1126), .ZN(n4225) );
  INV_X4 U7347 ( .A(n6954), .ZN(n6916) );
  OAI21_X2 U7348 ( .B1(n6634), .B2(n741), .A(n758), .ZN(n4226) );
  OAI21_X2 U7349 ( .B1(n6635), .B2(n373), .A(n390), .ZN(n4227) );
  OAI21_X2 U7350 ( .B1(n6634), .B2(n6760), .A(n289), .ZN(n4228) );
  INV_X4 U7351 ( .A(n6957), .ZN(n6936) );
  OAI21_X2 U7352 ( .B1(n6635), .B2(n237), .A(n254), .ZN(n4229) );
  OAI21_X2 U7353 ( .B1(n5663), .B2(n6767), .A(n221), .ZN(n4230) );
  OAI21_X2 U7354 ( .B1(n6634), .B2(n6770), .A(n187), .ZN(n4231) );
  OAI21_X2 U7355 ( .B1(n5663), .B2(n6774), .A(n152), .ZN(n4232) );
  OAI21_X2 U7356 ( .B1(n5663), .B2(n6777), .A(n118), .ZN(n4233) );
  OAI21_X2 U7357 ( .B1(n34), .B2(n5663), .A(n68), .ZN(n4234) );
  OAI21_X2 U7358 ( .B1(n6634), .B2(net367597), .A(n1093), .ZN(n4235) );
  OAI21_X2 U7359 ( .B1(n6634), .B2(n1043), .A(n1060), .ZN(n4236) );
  OAI21_X2 U7360 ( .B1(n6634), .B2(n6688), .A(n1026), .ZN(n4237) );
  OAI21_X2 U7361 ( .B1(n6634), .B2(n6691), .A(n992), .ZN(n4238) );
  INV_X4 U7362 ( .A(n6953), .ZN(n6908) );
  OAI21_X2 U7363 ( .B1(n6634), .B2(n942), .A(n959), .ZN(n4239) );
  OAI21_X2 U7364 ( .B1(n6634), .B2(n6702), .A(n891), .ZN(n4241) );
  OAI21_X2 U7365 ( .B1(n6634), .B2(n6706), .A(n858), .ZN(n4242) );
  OAI21_X2 U7366 ( .B1(n6634), .B2(n6712), .A(n791), .ZN(n4244) );
  OAI21_X2 U7367 ( .B1(n6635), .B2(n708), .A(n725), .ZN(n4245) );
  OAI21_X2 U7368 ( .B1(n6635), .B2(n675), .A(n692), .ZN(n4246) );
  INV_X4 U7369 ( .A(n6955), .ZN(n6924) );
  OAI21_X2 U7370 ( .B1(n6635), .B2(n540), .A(n557), .ZN(n4250) );
  INV_X4 U7371 ( .A(n6955), .ZN(n6928) );
  OAI21_X2 U7372 ( .B1(n6635), .B2(n439), .A(n456), .ZN(n4253) );
  OAI21_X2 U7373 ( .B1(n6635), .B2(n6751), .A(n423), .ZN(n4254) );
  OAI21_X2 U7374 ( .B1(n6632), .B2(n6679), .A(n1125), .ZN(n4258) );
  OAI21_X2 U7375 ( .B1(n6632), .B2(n6714), .A(n757), .ZN(n4259) );
  OAI21_X2 U7376 ( .B1(n6633), .B2(net367217), .A(n389), .ZN(n4260) );
  OAI21_X2 U7377 ( .B1(n6632), .B2(n6759), .A(n288), .ZN(n4261) );
  OAI21_X2 U7378 ( .B1(n5664), .B2(n6762), .A(n253), .ZN(n4262) );
  OAI21_X2 U7379 ( .B1(n6633), .B2(n6766), .A(n220), .ZN(n4263) );
  OAI21_X2 U7380 ( .B1(n5664), .B2(n6769), .A(n186), .ZN(n4264) );
  OAI21_X2 U7381 ( .B1(n6632), .B2(n6773), .A(n151), .ZN(n4265) );
  OAI21_X2 U7382 ( .B1(n5664), .B2(n6776), .A(n117), .ZN(n4266) );
  OAI21_X2 U7383 ( .B1(n6780), .B2(n5664), .A(n66), .ZN(n4267) );
  OAI21_X2 U7384 ( .B1(n6632), .B2(net367595), .A(n1092), .ZN(n4268) );
  OAI21_X2 U7385 ( .B1(n6632), .B2(n6684), .A(n1059), .ZN(n4269) );
  OAI21_X2 U7386 ( .B1(n6632), .B2(n6687), .A(n1025), .ZN(n4270) );
  OAI21_X2 U7387 ( .B1(n6632), .B2(n6690), .A(n991), .ZN(n4271) );
  OAI21_X2 U7388 ( .B1(n6632), .B2(n6694), .A(n958), .ZN(n4272) );
  OAI21_X2 U7389 ( .B1(n6632), .B2(n6698), .A(n924), .ZN(n4273) );
  OAI21_X2 U7390 ( .B1(n6632), .B2(n6701), .A(n890), .ZN(n4274) );
  OAI21_X2 U7391 ( .B1(n6632), .B2(n6705), .A(n857), .ZN(n4275) );
  OAI21_X2 U7392 ( .B1(n6632), .B2(n6708), .A(n824), .ZN(n4276) );
  OAI21_X2 U7393 ( .B1(n6632), .B2(n6711), .A(n790), .ZN(n4277) );
  OAI21_X2 U7394 ( .B1(n6633), .B2(n6718), .A(n724), .ZN(n4278) );
  OAI21_X2 U7395 ( .B1(n6633), .B2(n6723), .A(n691), .ZN(n4279) );
  OAI21_X2 U7396 ( .B1(n6633), .B2(n6726), .A(n658), .ZN(n4280) );
  OAI21_X2 U7397 ( .B1(n6633), .B2(n6729), .A(n624), .ZN(n4281) );
  OAI21_X2 U7398 ( .B1(n6633), .B2(n6733), .A(n589), .ZN(n4282) );
  OAI21_X2 U7399 ( .B1(n6633), .B2(n6737), .A(n556), .ZN(n4283) );
  OAI21_X2 U7400 ( .B1(n6633), .B2(n6741), .A(n523), .ZN(n4284) );
  OAI21_X2 U7401 ( .B1(n6633), .B2(n6744), .A(n489), .ZN(n4285) );
  OAI21_X2 U7402 ( .B1(n6633), .B2(n6747), .A(n455), .ZN(n4286) );
  OAI21_X2 U7403 ( .B1(n6633), .B2(n6750), .A(n422), .ZN(n4287) );
  OAI21_X2 U7404 ( .B1(n6633), .B2(n6753), .A(n356), .ZN(n4288) );
  OAI21_X2 U7405 ( .B1(n5664), .B2(n6756), .A(n322), .ZN(n4289) );
  AOI222_X1 U7406 ( .A1(n1147), .A2(drData[7]), .B1(daddr[7]), .B2(n1146), 
        .C1(aluJAL), .C2(aluPC8[7]), .ZN(n1232) );
  OAI21_X2 U7407 ( .B1(n6630), .B2(n6679), .A(n1124), .ZN(n4291) );
  OAI21_X2 U7408 ( .B1(n6630), .B2(n6714), .A(n756), .ZN(n4292) );
  OAI21_X2 U7409 ( .B1(n6631), .B2(net367217), .A(n388), .ZN(n4293) );
  OAI21_X2 U7410 ( .B1(n6631), .B2(n6759), .A(n287), .ZN(n4294) );
  OAI21_X2 U7411 ( .B1(n5665), .B2(n6762), .A(n252), .ZN(n4295) );
  OAI21_X2 U7412 ( .B1(n6630), .B2(n6766), .A(n219), .ZN(n4296) );
  OAI21_X2 U7413 ( .B1(n5665), .B2(n6769), .A(n185), .ZN(n4297) );
  OAI21_X2 U7414 ( .B1(n5665), .B2(n6773), .A(n150), .ZN(n4298) );
  OAI21_X2 U7415 ( .B1(n5665), .B2(n6776), .A(n116), .ZN(n4299) );
  OAI21_X2 U7416 ( .B1(n6780), .B2(n5665), .A(n64), .ZN(n4300) );
  OAI21_X2 U7417 ( .B1(n6630), .B2(net367595), .A(n1091), .ZN(n4301) );
  OAI21_X2 U7418 ( .B1(n6630), .B2(n6684), .A(n1058), .ZN(n4302) );
  OAI21_X2 U7419 ( .B1(n6630), .B2(n6687), .A(n1024), .ZN(n4303) );
  OAI21_X2 U7420 ( .B1(n6630), .B2(n6690), .A(n990), .ZN(n4304) );
  OAI21_X2 U7421 ( .B1(n6630), .B2(n6694), .A(n957), .ZN(n4305) );
  OAI21_X2 U7422 ( .B1(n6630), .B2(n6698), .A(n923), .ZN(n4306) );
  OAI21_X2 U7423 ( .B1(n6630), .B2(n6701), .A(n889), .ZN(n4307) );
  OAI21_X2 U7424 ( .B1(n6630), .B2(n6705), .A(n856), .ZN(n4308) );
  OAI21_X2 U7425 ( .B1(n6630), .B2(n6708), .A(n823), .ZN(n4309) );
  OAI21_X2 U7426 ( .B1(n6630), .B2(n6711), .A(n789), .ZN(n4310) );
  OAI21_X2 U7427 ( .B1(n6631), .B2(n6718), .A(n723), .ZN(n4311) );
  OAI21_X2 U7428 ( .B1(n6631), .B2(n6723), .A(n690), .ZN(n4312) );
  OAI21_X2 U7429 ( .B1(n6631), .B2(n6726), .A(n657), .ZN(n4313) );
  OAI21_X2 U7430 ( .B1(n6631), .B2(n6729), .A(n623), .ZN(n4314) );
  OAI21_X2 U7431 ( .B1(n6631), .B2(n6733), .A(n588), .ZN(n4315) );
  OAI21_X2 U7432 ( .B1(n6631), .B2(n6737), .A(n555), .ZN(n4316) );
  OAI21_X2 U7433 ( .B1(n6631), .B2(n6741), .A(n522), .ZN(n4317) );
  OAI21_X2 U7434 ( .B1(n6631), .B2(n6744), .A(n488), .ZN(n4318) );
  OAI21_X2 U7435 ( .B1(n6631), .B2(n6747), .A(n454), .ZN(n4319) );
  OAI21_X2 U7436 ( .B1(n6631), .B2(n6750), .A(n421), .ZN(n4320) );
  OAI21_X2 U7437 ( .B1(n6631), .B2(n6753), .A(n355), .ZN(n4321) );
  OAI21_X2 U7438 ( .B1(n6630), .B2(n6756), .A(n321), .ZN(n4322) );
  OAI21_X2 U7439 ( .B1(n5689), .B2(n5358), .A(n1234), .ZN(n4323) );
  OAI21_X2 U7440 ( .B1(n6628), .B2(n6679), .A(n1123), .ZN(n4324) );
  OAI21_X2 U7441 ( .B1(n6628), .B2(n6714), .A(n755), .ZN(n4325) );
  OAI21_X2 U7442 ( .B1(n6629), .B2(net367217), .A(n387), .ZN(n4326) );
  OAI21_X2 U7443 ( .B1(n5666), .B2(n6759), .A(n286), .ZN(n4327) );
  OAI21_X2 U7444 ( .B1(n5666), .B2(n6762), .A(n251), .ZN(n4328) );
  OAI21_X2 U7445 ( .B1(n5666), .B2(n6766), .A(n218), .ZN(n4329) );
  OAI21_X2 U7446 ( .B1(n6629), .B2(n6769), .A(n184), .ZN(n4330) );
  OAI21_X2 U7447 ( .B1(n5666), .B2(n6773), .A(n149), .ZN(n4331) );
  OAI21_X2 U7448 ( .B1(n6628), .B2(n6776), .A(n115), .ZN(n4332) );
  OAI21_X2 U7449 ( .B1(n6780), .B2(n5666), .A(n62), .ZN(n4333) );
  OAI21_X2 U7450 ( .B1(n6628), .B2(net367595), .A(n1090), .ZN(n4334) );
  OAI21_X2 U7451 ( .B1(n6628), .B2(n6684), .A(n1057), .ZN(n4335) );
  OAI21_X2 U7452 ( .B1(n6628), .B2(n6687), .A(n1023), .ZN(n4336) );
  OAI21_X2 U7453 ( .B1(n6628), .B2(n6690), .A(n989), .ZN(n4337) );
  OAI21_X2 U7454 ( .B1(n6628), .B2(n6694), .A(n956), .ZN(n4338) );
  OAI21_X2 U7455 ( .B1(n6628), .B2(n6701), .A(n888), .ZN(n4340) );
  INV_X4 U7456 ( .A(n6947), .ZN(n6862) );
  OAI21_X2 U7457 ( .B1(n6628), .B2(n6705), .A(n855), .ZN(n4341) );
  OAI21_X2 U7458 ( .B1(n6628), .B2(n6708), .A(n822), .ZN(n4342) );
  OAI21_X2 U7459 ( .B1(n6628), .B2(n6711), .A(n788), .ZN(n4343) );
  OAI21_X2 U7460 ( .B1(n6629), .B2(n6718), .A(n722), .ZN(n4344) );
  OAI21_X2 U7461 ( .B1(n6629), .B2(n6723), .A(n689), .ZN(n4345) );
  INV_X4 U7462 ( .A(n6946), .ZN(n6854) );
  OAI21_X2 U7463 ( .B1(n6629), .B2(n6726), .A(n656), .ZN(n4346) );
  OAI21_X2 U7464 ( .B1(n6629), .B2(n6729), .A(n622), .ZN(n4347) );
  OAI21_X2 U7465 ( .B1(n6629), .B2(n6733), .A(n587), .ZN(n4348) );
  OAI21_X2 U7466 ( .B1(n6629), .B2(n6737), .A(n554), .ZN(n4349) );
  OAI21_X2 U7467 ( .B1(n6629), .B2(n6741), .A(n521), .ZN(n4350) );
  OAI21_X2 U7468 ( .B1(n6629), .B2(n6744), .A(n487), .ZN(n4351) );
  OAI21_X2 U7469 ( .B1(n6629), .B2(n6747), .A(n453), .ZN(n4352) );
  OAI21_X2 U7470 ( .B1(n6629), .B2(n6750), .A(n420), .ZN(n4353) );
  OAI21_X2 U7471 ( .B1(n6629), .B2(n6753), .A(n354), .ZN(n4354) );
  OAI21_X2 U7472 ( .B1(n6628), .B2(n6756), .A(n320), .ZN(n4355) );
  OAI21_X2 U7473 ( .B1(n5689), .B2(n5357), .A(n1236), .ZN(n4356) );
  OAI21_X2 U7474 ( .B1(n6626), .B2(n6679), .A(n1122), .ZN(n4357) );
  OAI21_X2 U7475 ( .B1(n6626), .B2(n6714), .A(n754), .ZN(n4358) );
  OAI21_X2 U7476 ( .B1(n6627), .B2(net367217), .A(n386), .ZN(n4359) );
  OAI21_X2 U7477 ( .B1(n5667), .B2(n6759), .A(n285), .ZN(n4360) );
  OAI21_X2 U7478 ( .B1(n6626), .B2(n6762), .A(n250), .ZN(n4361) );
  OAI21_X2 U7479 ( .B1(n5667), .B2(n6766), .A(n217), .ZN(n4362) );
  OAI21_X2 U7480 ( .B1(n5667), .B2(n6769), .A(n183), .ZN(n4363) );
  OAI21_X2 U7481 ( .B1(n5667), .B2(n6773), .A(n148), .ZN(n4364) );
  OAI21_X2 U7482 ( .B1(n6626), .B2(n6776), .A(n114), .ZN(n4365) );
  OAI21_X2 U7483 ( .B1(n6780), .B2(n5667), .A(n60), .ZN(n4366) );
  OAI21_X2 U7484 ( .B1(n6626), .B2(net367595), .A(n1089), .ZN(n4367) );
  OAI21_X2 U7485 ( .B1(n6626), .B2(n6684), .A(n1056), .ZN(n4368) );
  OAI21_X2 U7486 ( .B1(n6626), .B2(n6687), .A(n1022), .ZN(n4369) );
  OAI21_X2 U7487 ( .B1(n6626), .B2(n6690), .A(n988), .ZN(n4370) );
  OAI21_X2 U7488 ( .B1(n6626), .B2(n6694), .A(n955), .ZN(n4371) );
  OAI21_X2 U7489 ( .B1(n6626), .B2(n6698), .A(n921), .ZN(n4372) );
  OAI21_X2 U7490 ( .B1(n6626), .B2(n6705), .A(n854), .ZN(n4374) );
  OAI21_X2 U7491 ( .B1(n6626), .B2(n6708), .A(n821), .ZN(n4375) );
  OAI21_X2 U7492 ( .B1(n6626), .B2(n6711), .A(n787), .ZN(n4376) );
  OAI21_X2 U7493 ( .B1(n6627), .B2(n6718), .A(n721), .ZN(n4377) );
  OAI21_X2 U7494 ( .B1(n6627), .B2(n6723), .A(n688), .ZN(n4378) );
  OAI21_X2 U7495 ( .B1(n6627), .B2(n6726), .A(n655), .ZN(n4379) );
  OAI21_X2 U7496 ( .B1(n6627), .B2(n6729), .A(n621), .ZN(n4380) );
  OAI21_X2 U7497 ( .B1(n6627), .B2(n6737), .A(n553), .ZN(n4382) );
  OAI21_X2 U7498 ( .B1(n6627), .B2(n6741), .A(n520), .ZN(n4383) );
  OAI21_X2 U7499 ( .B1(n6627), .B2(n6744), .A(n486), .ZN(n4384) );
  OAI21_X2 U7500 ( .B1(n6627), .B2(n6747), .A(n452), .ZN(n4385) );
  OAI21_X2 U7501 ( .B1(n6627), .B2(n6750), .A(n419), .ZN(n4386) );
  OAI21_X2 U7502 ( .B1(n6627), .B2(n6753), .A(n353), .ZN(n4387) );
  OAI21_X2 U7503 ( .B1(n6627), .B2(n6756), .A(n319), .ZN(n4388) );
  OAI21_X2 U7504 ( .B1(n5689), .B2(n5356), .A(n1238), .ZN(n4389) );
  OAI21_X2 U7505 ( .B1(n6624), .B2(n6679), .A(n1121), .ZN(n4390) );
  INV_X4 U7506 ( .A(n6956), .ZN(n6858) );
  OAI21_X2 U7507 ( .B1(n6624), .B2(n6714), .A(n753), .ZN(n4391) );
  OAI21_X2 U7508 ( .B1(n6625), .B2(net367217), .A(n385), .ZN(n4392) );
  OAI21_X2 U7509 ( .B1(n5668), .B2(n6759), .A(n284), .ZN(n4393) );
  OAI21_X2 U7510 ( .B1(n5668), .B2(n6762), .A(n249), .ZN(n4394) );
  OAI21_X2 U7511 ( .B1(n6625), .B2(n6766), .A(n216), .ZN(n4395) );
  OAI21_X2 U7512 ( .B1(n5668), .B2(n6769), .A(n182), .ZN(n4396) );
  OAI21_X2 U7513 ( .B1(n6624), .B2(n6773), .A(n147), .ZN(n4397) );
  OAI21_X2 U7514 ( .B1(n5668), .B2(n6776), .A(n113), .ZN(n4398) );
  OAI21_X2 U7515 ( .B1(n6780), .B2(n5668), .A(n58), .ZN(n4399) );
  INV_X4 U7516 ( .A(n6948), .ZN(n6870) );
  OAI21_X2 U7517 ( .B1(n6624), .B2(n6684), .A(n1055), .ZN(n4401) );
  OAI21_X2 U7518 ( .B1(n6624), .B2(n6687), .A(n1021), .ZN(n4402) );
  OAI21_X2 U7519 ( .B1(n6624), .B2(n6690), .A(n987), .ZN(n4403) );
  INV_X4 U7520 ( .A(n6948), .ZN(n6866) );
  OAI21_X2 U7521 ( .B1(n6624), .B2(n6694), .A(n954), .ZN(n4404) );
  OAI21_X2 U7522 ( .B1(n6624), .B2(n6698), .A(n920), .ZN(n4405) );
  OAI21_X2 U7523 ( .B1(n6624), .B2(n6701), .A(n886), .ZN(n4406) );
  OAI21_X2 U7524 ( .B1(n6625), .B2(n6718), .A(n720), .ZN(n4410) );
  OAI21_X2 U7525 ( .B1(n6625), .B2(n6723), .A(n687), .ZN(n4411) );
  OAI21_X2 U7526 ( .B1(n6625), .B2(n6729), .A(n620), .ZN(n4413) );
  OAI21_X2 U7527 ( .B1(n6625), .B2(n6737), .A(n552), .ZN(n4415) );
  OAI21_X2 U7528 ( .B1(n6625), .B2(n6744), .A(n485), .ZN(n4417) );
  INV_X4 U7529 ( .A(n6945), .ZN(n6846) );
  OAI21_X2 U7530 ( .B1(n6625), .B2(n6747), .A(n451), .ZN(n4418) );
  OAI21_X2 U7531 ( .B1(n6625), .B2(n6750), .A(n418), .ZN(n4419) );
  INV_X4 U7532 ( .A(n6950), .ZN(n6843) );
  OAI21_X2 U7533 ( .B1(n6625), .B2(n6753), .A(n352), .ZN(n4420) );
  OAI21_X2 U7534 ( .B1(n6625), .B2(n6756), .A(n318), .ZN(n4421) );
  OAI21_X2 U7535 ( .B1(n5689), .B2(n5362), .A(n1145), .ZN(n4422) );
  OAI21_X2 U7536 ( .B1(n6623), .B2(n6679), .A(n1120), .ZN(n4423) );
  OAI21_X2 U7537 ( .B1(n6623), .B2(n6714), .A(n752), .ZN(n4424) );
  OAI21_X2 U7538 ( .B1(n6623), .B2(net367217), .A(n384), .ZN(n4425) );
  OAI21_X2 U7539 ( .B1(n6623), .B2(n6759), .A(n283), .ZN(n4426) );
  OAI21_X2 U7540 ( .B1(n5682), .B2(n6762), .A(n248), .ZN(n4427) );
  OAI21_X2 U7541 ( .B1(n6623), .B2(n6766), .A(n215), .ZN(n4428) );
  OAI21_X2 U7542 ( .B1(n5682), .B2(n6773), .A(n146), .ZN(n4430) );
  OAI21_X2 U7543 ( .B1(n6623), .B2(n6776), .A(n112), .ZN(n4431) );
  OAI21_X2 U7544 ( .B1(n6780), .B2(n5682), .A(n56), .ZN(n4432) );
  OAI21_X2 U7545 ( .B1(n6623), .B2(net367595), .A(n1087), .ZN(n4433) );
  OAI21_X2 U7546 ( .B1(n6623), .B2(n6687), .A(n1020), .ZN(n4435) );
  OAI21_X2 U7547 ( .B1(n6623), .B2(n6690), .A(n986), .ZN(n4436) );
  OAI21_X2 U7548 ( .B1(n5682), .B2(n6698), .A(n919), .ZN(n4438) );
  OAI21_X2 U7549 ( .B1(n6623), .B2(n6701), .A(n885), .ZN(n4439) );
  OAI21_X2 U7550 ( .B1(n6623), .B2(n6705), .A(n852), .ZN(n4440) );
  OAI21_X2 U7551 ( .B1(n6623), .B2(n6708), .A(n819), .ZN(n4441) );
  OAI21_X2 U7552 ( .B1(n5682), .B2(n6711), .A(n785), .ZN(n4442) );
  OAI21_X2 U7553 ( .B1(n6623), .B2(n6718), .A(n719), .ZN(n4443) );
  OAI21_X2 U7554 ( .B1(n6623), .B2(n6723), .A(n686), .ZN(n4444) );
  OAI21_X2 U7555 ( .B1(n6623), .B2(n6726), .A(n653), .ZN(n4445) );
  OAI21_X2 U7556 ( .B1(n6623), .B2(n6729), .A(n619), .ZN(n4446) );
  OAI21_X2 U7557 ( .B1(n6623), .B2(n6733), .A(n584), .ZN(n4447) );
  OAI21_X2 U7558 ( .B1(n6623), .B2(n6737), .A(n551), .ZN(n4448) );
  OAI21_X2 U7559 ( .B1(n6623), .B2(n6744), .A(n484), .ZN(n4450) );
  OAI21_X2 U7560 ( .B1(n6623), .B2(n6747), .A(n450), .ZN(n4451) );
  OAI21_X2 U7561 ( .B1(n6623), .B2(n6750), .A(n417), .ZN(n4452) );
  OAI21_X2 U7562 ( .B1(n5682), .B2(n6756), .A(n317), .ZN(n4454) );
  OAI21_X2 U7563 ( .B1(n5689), .B2(n5361), .A(n1149), .ZN(n4455) );
  INV_X4 U7564 ( .A(n6951), .ZN(n6902) );
  OAI21_X2 U7565 ( .B1(n6621), .B2(n6679), .A(n1118), .ZN(n4456) );
  INV_X4 U7566 ( .A(n6956), .ZN(n6917) );
  OAI21_X2 U7567 ( .B1(n6621), .B2(n6714), .A(n750), .ZN(n4457) );
  INV_X4 U7568 ( .A(n6956), .ZN(n6931) );
  OAI21_X2 U7569 ( .B1(n6622), .B2(net367217), .A(n382), .ZN(n4458) );
  OAI21_X2 U7570 ( .B1(n6622), .B2(n6759), .A(n281), .ZN(n4459) );
  INV_X4 U7571 ( .A(n6958), .ZN(n6937) );
  OAI21_X2 U7572 ( .B1(n5670), .B2(n6762), .A(n246), .ZN(n4460) );
  INV_X4 U7573 ( .A(n6957), .ZN(n6938) );
  OAI21_X2 U7574 ( .B1(n6621), .B2(n6766), .A(n213), .ZN(n4461) );
  INV_X4 U7575 ( .A(n6958), .ZN(n6939) );
  OAI21_X2 U7576 ( .B1(n5670), .B2(n6769), .A(n179), .ZN(n4462) );
  OAI21_X2 U7577 ( .B1(n5670), .B2(n6773), .A(n144), .ZN(n4463) );
  INV_X4 U7578 ( .A(n6958), .ZN(n6942) );
  OAI21_X2 U7579 ( .B1(n5670), .B2(n6776), .A(n110), .ZN(n4464) );
  OAI21_X2 U7580 ( .B1(n6780), .B2(n5670), .A(n52), .ZN(n4465) );
  OAI21_X2 U7581 ( .B1(n6621), .B2(net367595), .A(n1085), .ZN(n4466) );
  OAI21_X2 U7582 ( .B1(n6621), .B2(n6684), .A(n1052), .ZN(n4467) );
  INV_X4 U7583 ( .A(n6952), .ZN(n6906) );
  OAI21_X2 U7584 ( .B1(n6621), .B2(n6687), .A(n1018), .ZN(n4468) );
  INV_X4 U7585 ( .A(n6952), .ZN(n6907) );
  OAI21_X2 U7586 ( .B1(n6621), .B2(n6690), .A(n984), .ZN(n4469) );
  INV_X4 U7587 ( .A(n6953), .ZN(n6909) );
  OAI21_X2 U7588 ( .B1(n6621), .B2(n6694), .A(n951), .ZN(n4470) );
  INV_X4 U7589 ( .A(n6953), .ZN(n6910) );
  OAI21_X2 U7590 ( .B1(n6621), .B2(n6698), .A(n917), .ZN(n4471) );
  OAI21_X2 U7591 ( .B1(n6621), .B2(n6701), .A(n883), .ZN(n4472) );
  INV_X4 U7592 ( .A(n6954), .ZN(n6913) );
  OAI21_X2 U7593 ( .B1(n6621), .B2(n6705), .A(n850), .ZN(n4473) );
  OAI21_X2 U7594 ( .B1(n6621), .B2(n6708), .A(n817), .ZN(n4474) );
  INV_X4 U7595 ( .A(n6954), .ZN(n6915) );
  OAI21_X2 U7596 ( .B1(n6621), .B2(n6711), .A(n783), .ZN(n4475) );
  INV_X4 U7597 ( .A(n6954), .ZN(n6918) );
  OAI21_X2 U7598 ( .B1(n6622), .B2(n6718), .A(n717), .ZN(n4476) );
  INV_X4 U7599 ( .A(n6954), .ZN(n6919) );
  OAI21_X2 U7600 ( .B1(n6622), .B2(n6723), .A(n684), .ZN(n4477) );
  OAI21_X2 U7601 ( .B1(n6622), .B2(n6726), .A(n651), .ZN(n4478) );
  INV_X4 U7602 ( .A(n6953), .ZN(n6922) );
  OAI21_X2 U7603 ( .B1(n6622), .B2(n6729), .A(n617), .ZN(n4479) );
  INV_X4 U7604 ( .A(n6955), .ZN(n6923) );
  OAI21_X2 U7605 ( .B1(n6622), .B2(n6733), .A(n582), .ZN(n4480) );
  INV_X4 U7606 ( .A(n6955), .ZN(n6925) );
  OAI21_X2 U7607 ( .B1(n6622), .B2(n6737), .A(n549), .ZN(n4481) );
  INV_X4 U7608 ( .A(n6955), .ZN(n6926) );
  OAI21_X2 U7609 ( .B1(n6622), .B2(n6741), .A(n516), .ZN(n4482) );
  OAI21_X2 U7610 ( .B1(n6622), .B2(n6744), .A(n482), .ZN(n4483) );
  OAI21_X2 U7611 ( .B1(n6622), .B2(n6747), .A(n448), .ZN(n4484) );
  INV_X4 U7612 ( .A(n6956), .ZN(n6930) );
  OAI21_X2 U7613 ( .B1(n6622), .B2(n6750), .A(n415), .ZN(n4485) );
  INV_X4 U7614 ( .A(n6957), .ZN(n6933) );
  OAI21_X2 U7615 ( .B1(n6622), .B2(n6753), .A(n349), .ZN(n4486) );
  INV_X4 U7616 ( .A(n6957), .ZN(n6934) );
  OAI21_X2 U7617 ( .B1(n6621), .B2(n6756), .A(n315), .ZN(n4487) );
  OAI21_X2 U7618 ( .B1(n5689), .B2(n5360), .A(n1151), .ZN(n4488) );
  INV_X4 U7619 ( .A(n6949), .ZN(n6872) );
  OAI21_X2 U7620 ( .B1(n6620), .B2(n6678), .A(n1117), .ZN(n4489) );
  OAI21_X2 U7621 ( .B1(n6620), .B2(n6713), .A(n749), .ZN(n4490) );
  OAI21_X2 U7622 ( .B1(n5683), .B2(n6758), .A(n280), .ZN(n4492) );
  OAI21_X2 U7623 ( .B1(n6620), .B2(n6761), .A(n245), .ZN(n4493) );
  INV_X4 U7624 ( .A(n6948), .ZN(n6837) );
  OAI21_X2 U7625 ( .B1(n5683), .B2(n6765), .A(n212), .ZN(n4494) );
  OAI21_X2 U7626 ( .B1(n6620), .B2(n6768), .A(n178), .ZN(n4495) );
  OAI21_X2 U7627 ( .B1(n5683), .B2(n6772), .A(n143), .ZN(n4496) );
  OAI21_X2 U7628 ( .B1(n6779), .B2(n5683), .A(n50), .ZN(n4498) );
  INV_X4 U7629 ( .A(n6948), .ZN(n6869) );
  OAI21_X2 U7630 ( .B1(n6620), .B2(n6683), .A(n1051), .ZN(n4500) );
  OAI21_X2 U7631 ( .B1(n5683), .B2(n6686), .A(n1017), .ZN(n4501) );
  OAI21_X2 U7632 ( .B1(n6620), .B2(n6689), .A(n983), .ZN(n4502) );
  OAI21_X2 U7633 ( .B1(n6620), .B2(n6693), .A(n950), .ZN(n4503) );
  OAI21_X2 U7634 ( .B1(n5683), .B2(n6697), .A(n916), .ZN(n4504) );
  INV_X4 U7635 ( .A(n6947), .ZN(n6863) );
  OAI21_X2 U7636 ( .B1(n6620), .B2(n6700), .A(n882), .ZN(n4505) );
  OAI21_X2 U7637 ( .B1(n6620), .B2(n6704), .A(n849), .ZN(n4506) );
  INV_X4 U7638 ( .A(n6954), .ZN(n6860) );
  OAI21_X2 U7639 ( .B1(n5683), .B2(n6707), .A(n816), .ZN(n4507) );
  OAI21_X2 U7640 ( .B1(n6620), .B2(n6710), .A(n782), .ZN(n4508) );
  INV_X4 U7641 ( .A(n6957), .ZN(n6856) );
  OAI21_X2 U7642 ( .B1(n6620), .B2(n6717), .A(n716), .ZN(n4509) );
  INV_X4 U7643 ( .A(n6958), .ZN(n6855) );
  OAI21_X2 U7644 ( .B1(n6620), .B2(n6722), .A(n683), .ZN(n4510) );
  INV_X4 U7645 ( .A(n6946), .ZN(n6853) );
  OAI21_X2 U7646 ( .B1(n6620), .B2(n6725), .A(n650), .ZN(n4511) );
  OAI21_X2 U7647 ( .B1(n6620), .B2(n6728), .A(n616), .ZN(n4512) );
  INV_X4 U7648 ( .A(n6946), .ZN(n6851) );
  OAI21_X2 U7649 ( .B1(n6620), .B2(n6732), .A(n581), .ZN(n4513) );
  OAI21_X2 U7650 ( .B1(n6620), .B2(n6736), .A(n548), .ZN(n4514) );
  OAI21_X2 U7651 ( .B1(n6620), .B2(n6740), .A(n515), .ZN(n4515) );
  OAI21_X2 U7652 ( .B1(n6620), .B2(n6743), .A(n481), .ZN(n4516) );
  OAI21_X2 U7653 ( .B1(n6620), .B2(n6748), .A(n447), .ZN(n4517) );
  OAI21_X2 U7654 ( .B1(n6620), .B2(n6749), .A(n414), .ZN(n4518) );
  OAI21_X2 U7655 ( .B1(n6620), .B2(n6752), .A(n348), .ZN(n4519) );
  OAI21_X2 U7656 ( .B1(n6620), .B2(n6755), .A(n314), .ZN(n4520) );
  OAI21_X2 U7657 ( .B1(n5689), .B2(n5359), .A(n1153), .ZN(n4521) );
  INV_X4 U7658 ( .A(n6949), .ZN(n6873) );
  INV_X4 U7659 ( .A(n6951), .ZN(n6901) );
  INV_X4 U7660 ( .A(n6949), .ZN(n6874) );
  OAI21_X2 U7661 ( .B1(n6601), .B2(n12610), .A(n12609), .ZN(n4557) );
  INV_X4 U7662 ( .A(n6954), .ZN(n6914) );
  INV_X4 U7663 ( .A(n6955), .ZN(n6859) );
  NOR2_X1 U7664 ( .A1(n5478), .A2(n12822), .ZN(n12817) );
  INV_X4 U7665 ( .A(n6956), .ZN(n6927) );
  AOI21_X1 U7666 ( .B1(ifOut_73_), .B2(n6593), .A(n12839), .ZN(n12836) );
  INV_X4 U7667 ( .A(n6951), .ZN(n6900) );
  AOI21_X2 U7668 ( .B1(ifOut_9_), .B2(n6593), .A(n12839), .ZN(n12844) );
  INV_X4 U7669 ( .A(n6949), .ZN(n6875) );
  INV_X4 U7670 ( .A(n6957), .ZN(n6935) );
  INV_X4 U7671 ( .A(n6951), .ZN(n6899) );
  INV_X4 U7672 ( .A(n6958), .ZN(n6941) );
  NAND3_X1 U7673 ( .A1(n6604), .A2(n12878), .A3(n12877), .ZN(n12880) );
  INV_X4 U7674 ( .A(n6946), .ZN(n6897) );
  INV_X4 U7675 ( .A(n6952), .ZN(n6877) );
  INV_X4 U7676 ( .A(n6951), .ZN(n6880) );
  INV_X4 U7677 ( .A(n6947), .ZN(n6842) );
  OAI21_X1 U7678 ( .B1(n12920), .B2(n13428), .A(n12919), .ZN(n4717) );
  OAI21_X1 U7679 ( .B1(ifInst[29]), .B2(n12917), .A(n13324), .ZN(n12918) );
  OAI21_X2 U7680 ( .B1(n12923), .B2(n13332), .A(n12922), .ZN(n4719) );
  NOR2_X2 U7681 ( .A1(n13497), .A2(n13322), .ZN(n12923) );
  INV_X4 U7682 ( .A(n6950), .ZN(n6886) );
  INV_X4 U7683 ( .A(n6947), .ZN(n6890) );
  NOR2_X2 U7684 ( .A1(n13249), .A2(net358618), .ZN(n13254) );
  INV_X4 U7685 ( .A(n6957), .ZN(n6883) );
  INV_X4 U7686 ( .A(n6948), .ZN(n6891) );
  INV_X4 U7687 ( .A(n6958), .ZN(n6940) );
  NAND3_X2 U7688 ( .A1(n13299), .A2(n13298), .A3(n13297), .ZN(n4782) );
  NAND3_X1 U7689 ( .A1(n13321), .A2(n13539), .A3(n13493), .ZN(n13328) );
  INV_X4 U7690 ( .A(n6956), .ZN(n6929) );
  NOR3_X2 U7691 ( .A1(n2082), .A2(ifInst[26]), .A3(n13358), .ZN(n13344) );
  NAND3_X2 U7692 ( .A1(n13355), .A2(n13354), .A3(n13353), .ZN(n4790) );
  INV_X4 U7693 ( .A(n6946), .ZN(n6852) );
  NAND3_X2 U7694 ( .A1(n13371), .A2(n13370), .A3(n13369), .ZN(n13608) );
  INV_X4 U7695 ( .A(n6950), .ZN(n6885) );
  INV_X4 U7696 ( .A(n6953), .ZN(n6889) );
  INV_X4 U7697 ( .A(n6954), .ZN(n6879) );
  NAND3_X1 U7698 ( .A1(ifInst[28]), .A2(n6581), .A3(n13396), .ZN(n13398) );
  NOR2_X2 U7699 ( .A1(n13403), .A2(n13402), .ZN(n4814) );
  NOR3_X1 U7700 ( .A1(ifInst[28]), .A2(n13539), .A3(n13400), .ZN(n13401) );
  INV_X4 U7701 ( .A(n6955), .ZN(n6881) );
  OAI21_X1 U7702 ( .B1(n13434), .B2(n5645), .A(n13406), .ZN(n4816) );
  INV_X4 U7703 ( .A(n6947), .ZN(n6861) );
  INV_X4 U7704 ( .A(n6947), .ZN(n6865) );
  INV_X4 U7705 ( .A(n6949), .ZN(n6892) );
  INV_X4 U7706 ( .A(n6956), .ZN(n6882) );
  NOR3_X1 U7707 ( .A1(n13434), .A2(n5455), .A3(n13427), .ZN(n4827) );
  INV_X4 U7708 ( .A(n6952), .ZN(n6893) );
  INV_X4 U7709 ( .A(n6951), .ZN(n6894) );
  INV_X4 U7710 ( .A(n6950), .ZN(n6895) );
  INV_X4 U7711 ( .A(n6949), .ZN(n6896) );
  INV_X4 U7712 ( .A(n6951), .ZN(n6876) );
  INV_X4 U7713 ( .A(n6951), .ZN(n6898) );
  INV_X4 U7714 ( .A(n6952), .ZN(n6921) );
  NOR2_X2 U7715 ( .A1(n5312), .A2(n13499), .ZN(n13500) );
  INV_X4 U7716 ( .A(n6958), .ZN(n6884) );
  INV_X4 U7717 ( .A(n6947), .ZN(n6864) );
  INV_X4 U7718 ( .A(n6948), .ZN(n6841) );
  INV_X4 U7719 ( .A(n6949), .ZN(n6871) );
  INV_X4 U7720 ( .A(n6952), .ZN(n6905) );
  INV_X4 U7721 ( .A(n6953), .ZN(n6878) );
  INV_X4 U7722 ( .A(n6953), .ZN(n6911) );
  INV_X4 U7723 ( .A(n6945), .ZN(n6849) );
  INV_X4 U7724 ( .A(n6945), .ZN(n6848) );
  INV_X4 U7725 ( .A(n6946), .ZN(n6845) );
  INV_X4 U7726 ( .A(n6952), .ZN(n6904) );
  INV_X4 U7727 ( .A(n6952), .ZN(n6903) );
  INV_X4 U7728 ( .A(n6953), .ZN(n6912) );
  INV_X4 U7729 ( .A(n6948), .ZN(n6868) );
  INV_X4 U7730 ( .A(n6948), .ZN(n6867) );
  INV_X4 U7731 ( .A(n6949), .ZN(n6836) );
  INV_X8 U7732 ( .A(n6816), .ZN(n6805) );
  INV_X4 U7733 ( .A(n6945), .ZN(n6840) );
  INV_X4 U7734 ( .A(n6945), .ZN(n6844) );
  INV_X4 U7735 ( .A(n6945), .ZN(n6847) );
  INV_X4 U7736 ( .A(regRst), .ZN(n6944) );
  INV_X4 U7737 ( .A(n6950), .ZN(n6888) );
  INV_X4 U7738 ( .A(n6950), .ZN(n6857) );
  INV_X4 U7739 ( .A(n6950), .ZN(n6887) );
  INV_X4 U7740 ( .A(net366967), .ZN(net375721) );
  INV_X8 U7741 ( .A(n6819), .ZN(n6815) );
  INV_X4 U7742 ( .A(regRst), .ZN(n6959) );
  INV_X4 U7743 ( .A(n6946), .ZN(n6839) );
  INV_X4 U7744 ( .A(n6946), .ZN(n6850) );
  INV_X4 U7745 ( .A(n6947), .ZN(n6838) );
  INV_X8 U7746 ( .A(n6817), .ZN(n6803) );
  INV_X4 U7747 ( .A(n6820), .ZN(n6819) );
  AND3_X4 U7748 ( .A1(idOut_22_), .A2(n9190), .A3(n9189), .ZN(n5288) );
  INV_X4 U7749 ( .A(n13231), .ZN(n6605) );
  AND2_X4 U7750 ( .A1(n203), .A2(n100), .ZN(n5289) );
  AND2_X4 U7751 ( .A1(n203), .A2(n169), .ZN(n5290) );
  INV_X4 U7752 ( .A(net366973), .ZN(net375547) );
  AND2_X4 U7753 ( .A1(n134), .A2(n100), .ZN(n5291) );
  AND2_X4 U7754 ( .A1(n807), .A2(n203), .ZN(n5292) );
  AND2_X4 U7755 ( .A1(n807), .A2(n168), .ZN(n5293) );
  AND2_X4 U7756 ( .A1(n641), .A2(n203), .ZN(n5294) );
  AND2_X4 U7757 ( .A1(n641), .A2(n168), .ZN(n5295) );
  AND2_X4 U7758 ( .A1(n506), .A2(n168), .ZN(n5296) );
  AND2_X4 U7759 ( .A1(n339), .A2(n168), .ZN(n5297) );
  AND2_X4 U7760 ( .A1(n305), .A2(n168), .ZN(n5298) );
  AND2_X4 U7761 ( .A1(n941), .A2(n134), .ZN(n5299) );
  AND2_X4 U7762 ( .A1(n941), .A2(n99), .ZN(n5300) );
  AND2_X4 U7763 ( .A1(n339), .A2(n99), .ZN(n5301) );
  AND2_X4 U7764 ( .A1(n807), .A2(n134), .ZN(n5302) );
  AND2_X4 U7765 ( .A1(n169), .A2(n99), .ZN(n5303) );
  INV_X2 U7766 ( .A(n13231), .ZN(n13062) );
  INV_X4 U7767 ( .A(n6560), .ZN(n6562) );
  INV_X4 U7768 ( .A(n5299), .ZN(n6688) );
  INV_X4 U7769 ( .A(n5300), .ZN(n6691) );
  INV_X4 U7770 ( .A(n5302), .ZN(n6702) );
  INV_X4 U7771 ( .A(n5303), .ZN(n6767) );
  INV_X4 U7772 ( .A(n5289), .ZN(net367597) );
  INV_X4 U7773 ( .A(n5290), .ZN(n6770) );
  INV_X4 U7774 ( .A(n5292), .ZN(n6709) );
  INV_X4 U7775 ( .A(n5298), .ZN(n6760) );
  INV_X4 U7776 ( .A(n5291), .ZN(n6777) );
  INV_X4 U7777 ( .A(n5294), .ZN(n6727) );
  INV_X4 U7778 ( .A(n5293), .ZN(n6712) );
  INV_X4 U7779 ( .A(n5301), .ZN(n6751) );
  INV_X4 U7780 ( .A(n5295), .ZN(n6730) );
  INV_X4 U7781 ( .A(n5297), .ZN(n6757) );
  INV_X4 U7782 ( .A(n5296), .ZN(n6745) );
  INV_X16 U7783 ( .A(n6828), .ZN(n6825) );
  INV_X16 U7784 ( .A(n6829), .ZN(n6823) );
  AND2_X4 U7785 ( .A1(n11520), .A2(n11519), .ZN(n5305) );
  INV_X4 U7786 ( .A(net369143), .ZN(n5770) );
  BUF_X4 U7787 ( .A(net369138), .Z(net369143) );
  AND2_X4 U7788 ( .A1(n12927), .A2(n6608), .ZN(n5306) );
  INV_X8 U7789 ( .A(n6600), .ZN(n6599) );
  INV_X8 U7790 ( .A(n6603), .ZN(n6602) );
  INV_X16 U7791 ( .A(n6603), .ZN(n6601) );
  INV_X16 U7792 ( .A(n6833), .ZN(n6832) );
  INV_X4 U7793 ( .A(net100619), .ZN(net367631) );
  INV_X4 U7794 ( .A(net366979), .ZN(net368862) );
  AND2_X2 U7795 ( .A1(n8710), .A2(n8709), .ZN(n5308) );
  INV_X4 U7796 ( .A(n13661), .ZN(n6608) );
  INV_X8 U7797 ( .A(n6608), .ZN(n6607) );
  INV_X4 U7798 ( .A(n5386), .ZN(n6560) );
  INV_X4 U7799 ( .A(regBoiz_N16), .ZN(n6820) );
  INV_X8 U7800 ( .A(n5331), .ZN(n6799) );
  INV_X4 U7801 ( .A(regRst), .ZN(n6946) );
  INV_X4 U7802 ( .A(regRst), .ZN(n6945) );
  NAND2_X4 U7803 ( .A1(n11726), .A2(n11727), .ZN(n5309) );
  NAND2_X4 U7804 ( .A1(n5821), .A2(net364941), .ZN(n5310) );
  OR2_X4 U7805 ( .A1(net375393), .A2(net364941), .ZN(n5311) );
  INV_X4 U7806 ( .A(n5354), .ZN(ifInst[25]) );
  AND2_X4 U7807 ( .A1(n12940), .A2(n6605), .ZN(n5315) );
  AND2_X4 U7808 ( .A1(idOut_25_), .A2(n6608), .ZN(n5316) );
  AND2_X4 U7809 ( .A1(n8706), .A2(n8705), .ZN(n5317) );
  INV_X4 U7810 ( .A(n6599), .ZN(n6604) );
  INV_X16 U7811 ( .A(n6833), .ZN(n6831) );
  INV_X16 U7812 ( .A(net368466), .ZN(net368467) );
  INV_X8 U7813 ( .A(regBoiz_N17), .ZN(n6828) );
  INV_X16 U7814 ( .A(n5389), .ZN(n6824) );
  INV_X4 U7815 ( .A(net359877), .ZN(net368205) );
  NAND2_X2 U7816 ( .A1(n6605), .A2(n13220), .ZN(n6554) );
  INV_X2 U7817 ( .A(n10043), .ZN(n6570) );
  INV_X4 U7818 ( .A(n6820), .ZN(n6818) );
  INV_X2 U7819 ( .A(n6819), .ZN(n6816) );
  INV_X4 U7820 ( .A(regRst), .ZN(n6950) );
  INV_X4 U7821 ( .A(regRst), .ZN(n6949) );
  INV_X4 U7822 ( .A(regRst), .ZN(n6948) );
  INV_X4 U7823 ( .A(regRst), .ZN(n6947) );
  AND2_X4 U7824 ( .A1(n10999), .A2(n13533), .ZN(n5332) );
  AND2_X4 U7825 ( .A1(net366987), .A2(n6795), .ZN(n5333) );
  AND2_X4 U7826 ( .A1(net377373), .A2(n11082), .ZN(n5334) );
  AND2_X2 U7827 ( .A1(n5573), .A2(net360919), .ZN(n5335) );
  AND2_X4 U7828 ( .A1(n12840), .A2(iaddr[2]), .ZN(n5347) );
  AND2_X4 U7829 ( .A1(ifOut_91_), .A2(ifInst[25]), .ZN(n5351) );
  XOR2_X2 U7830 ( .A(ifOut_88_), .B(ifInst[24]), .Z(n5352) );
  INV_X4 U7831 ( .A(n6610), .ZN(n6611) );
  INV_X4 U7832 ( .A(n13675), .ZN(n6609) );
  INV_X8 U7833 ( .A(n6591), .ZN(n6587) );
  NAND3_X2 U7834 ( .A1(n6608), .A2(n5314), .A3(n12939), .ZN(n13231) );
  AND2_X2 U7835 ( .A1(n13295), .A2(ifInst[28]), .ZN(n5380) );
  AND3_X4 U7836 ( .A1(n9196), .A2(n5345), .A3(n9677), .ZN(n5381) );
  AND2_X2 U7837 ( .A1(iaddr[6]), .A2(n12875), .ZN(n5385) );
  INV_X4 U7838 ( .A(net366919), .ZN(net376387) );
  AND2_X2 U7839 ( .A1(n9722), .A2(n9677), .ZN(n5386) );
  INV_X16 U7840 ( .A(net368571), .ZN(net368572) );
  NAND2_X2 U7841 ( .A1(n6605), .A2(n13220), .ZN(n6555) );
  NAND3_X2 U7842 ( .A1(didMult), .A2(n6608), .A3(n12945), .ZN(n5387) );
  AND2_X4 U7843 ( .A1(aluBoi_multOut[0]), .A2(n5690), .ZN(n5388) );
  INV_X4 U7844 ( .A(net367029), .ZN(net375614) );
  INV_X4 U7845 ( .A(regBoiz_N17), .ZN(n6829) );
  OR2_X4 U7846 ( .A1(n6549), .A2(n6571), .ZN(n5390) );
  NAND3_X1 U7847 ( .A1(n12926), .A2(n6608), .A3(n12925), .ZN(n13375) );
  INV_X4 U7848 ( .A(net368205), .ZN(net368203) );
  INV_X16 U7849 ( .A(net368203), .ZN(net368201) );
  NOR2_X2 U7850 ( .A1(n5519), .A2(aluJAL), .ZN(n1147) );
  INV_X4 U7851 ( .A(n10286), .ZN(n6572) );
  INV_X8 U7852 ( .A(n6572), .ZN(n6571) );
  INV_X4 U7853 ( .A(n5288), .ZN(n6563) );
  INV_X4 U7854 ( .A(n5288), .ZN(n6564) );
  INV_X4 U7855 ( .A(n6786), .ZN(n6230) );
  INV_X4 U7856 ( .A(n6786), .ZN(n6221) );
  INV_X4 U7857 ( .A(n1043), .ZN(n6682) );
  INV_X4 U7858 ( .A(n135), .ZN(n6771) );
  INV_X4 U7859 ( .A(n34), .ZN(n6778) );
  INV_X4 U7860 ( .A(n942), .ZN(n6692) );
  INV_X4 U7861 ( .A(n908), .ZN(n6696) );
  INV_X4 U7862 ( .A(n507), .ZN(n6739) );
  INV_X4 U7863 ( .A(n373), .ZN(net367231) );
  INV_X4 U7864 ( .A(n841), .ZN(n6703) );
  INV_X4 U7865 ( .A(n675), .ZN(n6721) );
  INV_X4 U7866 ( .A(n573), .ZN(n6731) );
  INV_X4 U7867 ( .A(n540), .ZN(n6735) );
  INV_X4 U7868 ( .A(n439), .ZN(n6746) );
  INV_X4 U7869 ( .A(net100619), .ZN(net368481) );
  XOR2_X1 U7870 ( .A(n5766), .B(n5768), .Z(n5392) );
  OR2_X4 U7871 ( .A1(aluBoi_aluBoi_shft_sraout[19]), .A2(
        aluBoi_aluBoi_shft_sraout[18]), .ZN(n5393) );
  INV_X4 U7872 ( .A(regRst), .ZN(n6954) );
  INV_X4 U7873 ( .A(regRst), .ZN(n6953) );
  INV_X4 U7874 ( .A(regRst), .ZN(n6952) );
  INV_X4 U7875 ( .A(regRst), .ZN(n6951) );
  OR2_X4 U7876 ( .A1(aluBoi_aluBoi_shft_sllout[21]), .A2(
        aluBoi_aluBoi_shft_sllout[20]), .ZN(n5394) );
  INV_X16 U7877 ( .A(n6510), .ZN(n6511) );
  INV_X2 U7878 ( .A(n6511), .ZN(n12060) );
  INV_X4 U7879 ( .A(n11258), .ZN(n11212) );
  XOR2_X2 U7880 ( .A(n10595), .B(n10593), .Z(n5395) );
  INV_X4 U7881 ( .A(n11231), .ZN(n10723) );
  INV_X4 U7882 ( .A(n5970), .ZN(n10941) );
  INV_X4 U7883 ( .A(net362050), .ZN(net362216) );
  INV_X4 U7884 ( .A(n12094), .ZN(n12086) );
  INV_X4 U7885 ( .A(n5884), .ZN(n11920) );
  XOR2_X2 U7886 ( .A(n11883), .B(n11882), .Z(n5403) );
  OR2_X2 U7887 ( .A1(n7942), .A2(n7941), .ZN(n5421) );
  OR2_X4 U7888 ( .A1(n7971), .A2(n7970), .ZN(n5422) );
  INV_X4 U7889 ( .A(n11124), .ZN(n11120) );
  AND2_X4 U7890 ( .A1(regBoiz_regfile_12__15_), .A2(net366919), .ZN(n5427) );
  AND2_X4 U7891 ( .A1(regBoiz_regfile_20__15_), .A2(net378321), .ZN(n5428) );
  AND2_X4 U7892 ( .A1(regBoiz_regfile_22__15_), .A2(net378321), .ZN(n5429) );
  AND2_X4 U7893 ( .A1(regBoiz_regfile_28__15_), .A2(net366919), .ZN(n5430) );
  AND2_X4 U7894 ( .A1(regBoiz_regfile_30__15_), .A2(net366933), .ZN(n5431) );
  AND2_X4 U7895 ( .A1(regBoiz_regfile_5__15_), .A2(net366933), .ZN(n5432) );
  AND2_X4 U7896 ( .A1(regBoiz_regfile_15__15_), .A2(net366919), .ZN(n5433) );
  AND2_X4 U7897 ( .A1(regBoiz_regfile_21__15_), .A2(net366933), .ZN(n5434) );
  AND2_X4 U7898 ( .A1(regBoiz_regfile_23__15_), .A2(net366939), .ZN(n5435) );
  AND2_X4 U7899 ( .A1(regBoiz_regfile_29__15_), .A2(net366939), .ZN(n5436) );
  AND2_X4 U7900 ( .A1(regBoiz_regfile_31__15_), .A2(net366939), .ZN(n5437) );
  AND2_X2 U7901 ( .A1(n6432), .A2(n11049), .ZN(n5438) );
  AND2_X4 U7902 ( .A1(n6241), .A2(n6242), .ZN(n5439) );
  OR2_X2 U7903 ( .A1(n8031), .A2(net366965), .ZN(n5440) );
  OR2_X4 U7904 ( .A1(net366967), .A2(n7976), .ZN(n5441) );
  AND2_X2 U7905 ( .A1(n11049), .A2(n11042), .ZN(n5442) );
  OR2_X4 U7906 ( .A1(n7990), .A2(net366965), .ZN(n5444) );
  OR2_X2 U7907 ( .A1(n7856), .A2(net366921), .ZN(n5445) );
  NAND2_X2 U7908 ( .A1(n12005), .A2(n12272), .ZN(n12021) );
  INV_X4 U7909 ( .A(net361312), .ZN(net361709) );
  AND2_X4 U7910 ( .A1(n7557), .A2(net366953), .ZN(n5446) );
  INV_X4 U7911 ( .A(n12289), .ZN(n12130) );
  AND2_X2 U7912 ( .A1(regBoiz_regfile_14__14_), .A2(net366939), .ZN(n5447) );
  AND2_X2 U7913 ( .A1(regBoiz_regfile_30__14_), .A2(net366939), .ZN(n5448) );
  AND3_X4 U7914 ( .A1(n9846), .A2(net367041), .A3(n9869), .ZN(n5449) );
  AND2_X2 U7915 ( .A1(regBoiz_regfile_14__15_), .A2(net366919), .ZN(n5450) );
  AND2_X2 U7916 ( .A1(regBoiz_regfile_28__21_), .A2(net366939), .ZN(n5451) );
  AND2_X2 U7917 ( .A1(regBoiz_regfile_30__21_), .A2(net366939), .ZN(n5452) );
  INV_X2 U7918 ( .A(n6423), .ZN(n6119) );
  OR2_X2 U7919 ( .A1(n7857), .A2(n5445), .ZN(n5453) );
  OR2_X2 U7920 ( .A1(n7981), .A2(n5440), .ZN(n5454) );
  INV_X4 U7921 ( .A(n12390), .ZN(n12558) );
  OR2_X4 U7922 ( .A1(n10043), .A2(n8834), .ZN(n5457) );
  AND2_X4 U7923 ( .A1(n12944), .A2(n6605), .ZN(n5460) );
  AND3_X4 U7924 ( .A1(ifInst[29]), .A2(n13422), .A3(n13325), .ZN(n5474) );
  AND2_X2 U7925 ( .A1(n13363), .A2(n5285), .ZN(n5492) );
  INV_X4 U7926 ( .A(n11787), .ZN(n5894) );
  INV_X4 U7927 ( .A(n11641), .ZN(n11644) );
  INV_X1 U7928 ( .A(n6548), .ZN(n6549) );
  INV_X4 U7929 ( .A(n10406), .ZN(n6577) );
  INV_X16 U7930 ( .A(n6577), .ZN(n6576) );
  AND2_X2 U7931 ( .A1(n7557), .A2(net378321), .ZN(n5553) );
  INV_X8 U7932 ( .A(n13430), .ZN(n6586) );
  AND3_X4 U7933 ( .A1(n5380), .A2(ifInst[26]), .A3(n13491), .ZN(n5555) );
  AND2_X4 U7934 ( .A1(ifOut_94_), .A2(n13488), .ZN(n5557) );
  INV_X8 U7935 ( .A(net368183), .ZN(net368181) );
  OR3_X1 U7936 ( .A1(ifInst[11]), .A2(ifInst[13]), .A3(ifInst[12]), .ZN(n5561)
         );
  OR2_X4 U7937 ( .A1(n2054), .A2(n13427), .ZN(n5575) );
  AND3_X4 U7938 ( .A1(n13221), .A2(n5927), .A3(n13220), .ZN(n5579) );
  INV_X8 U7939 ( .A(n5344), .ZN(n6835) );
  AND2_X2 U7940 ( .A1(regBoiz_regfile_29__31_), .A2(n6789), .ZN(n5586) );
  AND2_X2 U7941 ( .A1(regBoiz_regfile_31__31_), .A2(n6788), .ZN(n5587) );
  INV_X4 U7942 ( .A(n9677), .ZN(n5762) );
  AND2_X4 U7943 ( .A1(regBoiz_regfile_4__15_), .A2(net366939), .ZN(n5640) );
  AND2_X4 U7944 ( .A1(regBoiz_regfile_6__15_), .A2(net366939), .ZN(n5641) );
  NAND2_X2 U7945 ( .A1(n6605), .A2(n13220), .ZN(n13514) );
  INV_X4 U7946 ( .A(n13675), .ZN(n6610) );
  AND2_X4 U7947 ( .A1(regBoiz_regfile_7__15_), .A2(net366939), .ZN(n5642) );
  AND2_X4 U7948 ( .A1(regBoiz_regfile_13__15_), .A2(net378321), .ZN(n5643) );
  AND2_X2 U7949 ( .A1(regBoiz_regfile_7__21_), .A2(net366939), .ZN(n5644) );
  OR2_X4 U7950 ( .A1(n13539), .A2(n13427), .ZN(n5645) );
  NOR2_X2 U7951 ( .A1(aluJAL), .A2(aluMem2Reg), .ZN(n1146) );
  INV_X4 U7952 ( .A(wbBusWh[31]), .ZN(n6676) );
  INV_X4 U7953 ( .A(wbBusWh[31]), .ZN(n6677) );
  INV_X4 U7954 ( .A(wbBusWh[21]), .ZN(n6658) );
  INV_X4 U7955 ( .A(wbBusWh[20]), .ZN(n6656) );
  INV_X4 U7956 ( .A(wbBusWh[20]), .ZN(n6657) );
  INV_X4 U7957 ( .A(wbBusWh[19]), .ZN(n6655) );
  INV_X4 U7958 ( .A(wbBusWh[18]), .ZN(n6653) );
  INV_X4 U7959 ( .A(wbBusWh[18]), .ZN(n6654) );
  INV_X4 U7960 ( .A(wbBusWh[17]), .ZN(n6651) );
  INV_X4 U7961 ( .A(wbBusWh[17]), .ZN(n6652) );
  INV_X4 U7962 ( .A(wbBusWh[16]), .ZN(n6649) );
  INV_X4 U7963 ( .A(wbBusWh[16]), .ZN(n6650) );
  INV_X4 U7964 ( .A(wbBusWh[15]), .ZN(n6648) );
  INV_X4 U7965 ( .A(wbBusWh[15]), .ZN(n6647) );
  INV_X4 U7966 ( .A(wbBusWh[14]), .ZN(n6645) );
  INV_X4 U7967 ( .A(wbBusWh[14]), .ZN(n6646) );
  INV_X4 U7968 ( .A(wbBusWh[13]), .ZN(n6644) );
  INV_X4 U7969 ( .A(wbBusWh[12]), .ZN(n6642) );
  INV_X4 U7970 ( .A(wbBusWh[12]), .ZN(n6643) );
  INV_X4 U7971 ( .A(wbBusWh[30]), .ZN(n6674) );
  INV_X4 U7972 ( .A(wbBusWh[30]), .ZN(n6675) );
  INV_X4 U7973 ( .A(wbBusWh[11]), .ZN(n6640) );
  INV_X4 U7974 ( .A(wbBusWh[11]), .ZN(n6641) );
  INV_X4 U7975 ( .A(wbBusWh[10]), .ZN(n6638) );
  INV_X4 U7976 ( .A(wbBusWh[10]), .ZN(n6639) );
  INV_X4 U7977 ( .A(wbBusWh[9]), .ZN(n6637) );
  INV_X4 U7978 ( .A(wbBusWh[9]), .ZN(n6636) );
  INV_X4 U7979 ( .A(wbBusWh[8]), .ZN(n6634) );
  INV_X4 U7980 ( .A(wbBusWh[8]), .ZN(n6635) );
  INV_X4 U7981 ( .A(wbBusWh[7]), .ZN(n6632) );
  INV_X4 U7982 ( .A(wbBusWh[7]), .ZN(n6633) );
  INV_X4 U7983 ( .A(wbBusWh[6]), .ZN(n6630) );
  INV_X4 U7984 ( .A(wbBusWh[6]), .ZN(n6631) );
  INV_X4 U7985 ( .A(wbBusWh[5]), .ZN(n6628) );
  INV_X4 U7986 ( .A(wbBusWh[5]), .ZN(n6629) );
  INV_X4 U7987 ( .A(wbBusWh[4]), .ZN(n6626) );
  INV_X4 U7988 ( .A(wbBusWh[4]), .ZN(n6627) );
  INV_X4 U7989 ( .A(wbBusWh[3]), .ZN(n6625) );
  INV_X4 U7990 ( .A(wbBusWh[3]), .ZN(n6624) );
  INV_X4 U7991 ( .A(wbBusWh[29]), .ZN(n6672) );
  INV_X4 U7992 ( .A(wbBusWh[29]), .ZN(n6673) );
  INV_X4 U7993 ( .A(wbBusWh[1]), .ZN(n6621) );
  INV_X4 U7994 ( .A(wbBusWh[1]), .ZN(n6622) );
  INV_X4 U7995 ( .A(wbBusWh[28]), .ZN(n6670) );
  INV_X4 U7996 ( .A(wbBusWh[28]), .ZN(n6671) );
  INV_X4 U7997 ( .A(wbBusWh[26]), .ZN(n6666) );
  INV_X4 U7998 ( .A(wbBusWh[26]), .ZN(n6667) );
  INV_X4 U7999 ( .A(wbBusWh[24]), .ZN(n6663) );
  INV_X4 U8000 ( .A(wbBusWh[24]), .ZN(n6662) );
  INV_X4 U8001 ( .A(wbBusWh[23]), .ZN(n6661) );
  INV_X4 U8002 ( .A(wbBusWh[23]), .ZN(n6660) );
  INV_X4 U8003 ( .A(wbBusWh[22]), .ZN(n6659) );
  NAND3_X2 U8004 ( .A1(iaddr[11]), .A2(iaddr[10]), .A3(n12600), .ZN(n12816) );
  INV_X8 U8005 ( .A(regBoiz_N18), .ZN(n6833) );
  INV_X4 U8006 ( .A(wbBusWh[2]), .ZN(n6623) );
  INV_X4 U8007 ( .A(wbBusWh[0]), .ZN(n6620) );
  INV_X4 U8008 ( .A(wbBusWh[25]), .ZN(n6665) );
  INV_X4 U8009 ( .A(wbBusWh[25]), .ZN(n6664) );
  INV_X8 U8010 ( .A(net368518), .ZN(net368519) );
  INV_X1 U8011 ( .A(net368519), .ZN(net361631) );
  OR2_X4 U8012 ( .A1(n6569), .A2(n5462), .ZN(n5686) );
  INV_X4 U8013 ( .A(wbBusWh[27]), .ZN(n6668) );
  INV_X4 U8014 ( .A(wbBusWh[27]), .ZN(n6669) );
  NAND2_X1 U8015 ( .A1(n10331), .A2(iaddr[6]), .ZN(n12853) );
  INV_X4 U8016 ( .A(n5386), .ZN(n6561) );
  INV_X4 U8017 ( .A(n5387), .ZN(net368069) );
  AND2_X2 U8018 ( .A1(regBoiz_regfile_12__21_), .A2(net378321), .ZN(n5692) );
  AND2_X2 U8019 ( .A1(regBoiz_regfile_6__21_), .A2(net366939), .ZN(n5693) );
  AND2_X2 U8020 ( .A1(regBoiz_regfile_5__21_), .A2(net366919), .ZN(n5694) );
  AND2_X2 U8021 ( .A1(regBoiz_regfile_15__21_), .A2(net366919), .ZN(n5695) );
  INV_X4 U8022 ( .A(n13375), .ZN(n6579) );
  INV_X4 U8023 ( .A(n6579), .ZN(n6578) );
  INV_X16 U8024 ( .A(n6508), .ZN(n6509) );
  OR2_X4 U8025 ( .A1(n6569), .A2(n5512), .ZN(n5696) );
  INV_X4 U8026 ( .A(n13508), .ZN(n6600) );
  INV_X16 U8027 ( .A(n6530), .ZN(n6531) );
  INV_X2 U8028 ( .A(n6531), .ZN(n9822) );
  AND2_X2 U8029 ( .A1(regBoiz_regfile_20__21_), .A2(net366939), .ZN(n5697) );
  AND2_X2 U8030 ( .A1(regBoiz_regfile_21__21_), .A2(net378321), .ZN(n5698) );
  AND2_X2 U8031 ( .A1(regBoiz_regfile_29__21_), .A2(net366939), .ZN(n5699) );
  OR2_X4 U8032 ( .A1(n13309), .A2(n13408), .ZN(n5700) );
  INV_X4 U8033 ( .A(n5381), .ZN(n6567) );
  INV_X4 U8034 ( .A(n6567), .ZN(n6566) );
  OR2_X4 U8035 ( .A1(n11316), .A2(n6574), .ZN(n5701) );
  INV_X4 U8036 ( .A(net368445), .ZN(net368447) );
  INV_X4 U8037 ( .A(net368445), .ZN(net368446) );
  INV_X16 U8038 ( .A(n6550), .ZN(n6551) );
  INV_X16 U8039 ( .A(n6551), .ZN(n10369) );
  INV_X8 U8040 ( .A(net359750), .ZN(net368191) );
  INV_X8 U8041 ( .A(net368191), .ZN(net368185) );
  OR2_X2 U8042 ( .A1(n10372), .A2(n6574), .ZN(n5702) );
  INV_X16 U8043 ( .A(n6799), .ZN(n6814) );
  OR2_X4 U8044 ( .A1(n10346), .A2(n6574), .ZN(n5703) );
  INV_X16 U8045 ( .A(net369149), .ZN(net369240) );
  OR2_X4 U8046 ( .A1(n10189), .A2(n6574), .ZN(n5704) );
  OR2_X4 U8047 ( .A1(n11191), .A2(n6574), .ZN(n5705) );
  OR2_X4 U8048 ( .A1(n11003), .A2(n6574), .ZN(n5706) );
  OR2_X4 U8049 ( .A1(n10892), .A2(n6574), .ZN(n5707) );
  OR2_X4 U8050 ( .A1(n10708), .A2(n6574), .ZN(n5708) );
  OR2_X4 U8051 ( .A1(n10575), .A2(n6574), .ZN(n5709) );
  OR2_X4 U8052 ( .A1(n11380), .A2(n6573), .ZN(n5710) );
  OR2_X2 U8053 ( .A1(net361801), .A2(n6574), .ZN(n5711) );
  OR2_X2 U8054 ( .A1(n9729), .A2(n6573), .ZN(n5712) );
  OR2_X4 U8055 ( .A1(n9661), .A2(n9660), .ZN(n5713) );
  INV_X4 U8056 ( .A(n1109), .ZN(n6681) );
  INV_X4 U8057 ( .A(n6681), .ZN(n6678) );
  INV_X4 U8058 ( .A(n6681), .ZN(n6679) );
  INV_X4 U8059 ( .A(n6681), .ZN(n6680) );
  INV_X4 U8060 ( .A(n6682), .ZN(n6683) );
  INV_X4 U8061 ( .A(n6682), .ZN(n6684) );
  INV_X4 U8062 ( .A(n6682), .ZN(n6685) );
  INV_X4 U8063 ( .A(n5299), .ZN(n6686) );
  INV_X4 U8064 ( .A(n5299), .ZN(n6687) );
  INV_X4 U8065 ( .A(n5302), .ZN(n6701) );
  INV_X4 U8066 ( .A(n5302), .ZN(n6700) );
  INV_X4 U8067 ( .A(n5292), .ZN(n6708) );
  INV_X4 U8068 ( .A(n5292), .ZN(n6707) );
  INV_X4 U8069 ( .A(n5293), .ZN(n6711) );
  INV_X4 U8070 ( .A(n5293), .ZN(n6710) );
  INV_X4 U8071 ( .A(n741), .ZN(n6716) );
  INV_X4 U8072 ( .A(n6716), .ZN(n6713) );
  INV_X4 U8073 ( .A(n6716), .ZN(n6714) );
  INV_X4 U8074 ( .A(n6716), .ZN(n6715) );
  INV_X4 U8075 ( .A(n708), .ZN(n6720) );
  INV_X4 U8076 ( .A(n6720), .ZN(n6717) );
  INV_X4 U8077 ( .A(n6720), .ZN(n6718) );
  INV_X4 U8078 ( .A(n6720), .ZN(n6719) );
  INV_X4 U8079 ( .A(n6721), .ZN(n6722) );
  INV_X4 U8080 ( .A(n6721), .ZN(n6723) );
  INV_X4 U8081 ( .A(n6721), .ZN(n6724) );
  INV_X4 U8082 ( .A(n5294), .ZN(n6725) );
  INV_X4 U8083 ( .A(n5294), .ZN(n6726) );
  INV_X4 U8084 ( .A(n5295), .ZN(n6728) );
  INV_X4 U8085 ( .A(n5295), .ZN(n6729) );
  INV_X4 U8086 ( .A(n6731), .ZN(n6733) );
  INV_X4 U8087 ( .A(n6731), .ZN(n6732) );
  INV_X4 U8088 ( .A(n6731), .ZN(n6734) );
  INV_X4 U8089 ( .A(n5296), .ZN(n6743) );
  INV_X4 U8090 ( .A(n5296), .ZN(n6744) );
  INV_X4 U8091 ( .A(n5301), .ZN(n6749) );
  INV_X4 U8092 ( .A(n5301), .ZN(n6750) );
  INV_X4 U8093 ( .A(net367231), .ZN(net367215) );
  INV_X4 U8094 ( .A(net367231), .ZN(net367217) );
  INV_X4 U8095 ( .A(net367231), .ZN(net367221) );
  INV_X4 U8096 ( .A(n237), .ZN(n6764) );
  INV_X4 U8097 ( .A(n6764), .ZN(n6761) );
  INV_X4 U8098 ( .A(n6764), .ZN(n6762) );
  INV_X4 U8099 ( .A(n6764), .ZN(n6763) );
  INV_X4 U8100 ( .A(n5303), .ZN(n6765) );
  INV_X4 U8101 ( .A(n5303), .ZN(n6766) );
  INV_X4 U8102 ( .A(n5291), .ZN(n6775) );
  INV_X4 U8103 ( .A(n5291), .ZN(n6776) );
  INV_X4 U8104 ( .A(n6778), .ZN(n6779) );
  INV_X4 U8105 ( .A(n6778), .ZN(n6780) );
  INV_X4 U8106 ( .A(n6778), .ZN(n6781) );
  INV_X4 U8107 ( .A(n5289), .ZN(net367593) );
  INV_X4 U8108 ( .A(n5289), .ZN(net367595) );
  INV_X4 U8109 ( .A(n6703), .ZN(n6704) );
  INV_X4 U8110 ( .A(n6703), .ZN(n6705) );
  INV_X4 U8111 ( .A(n6703), .ZN(n6706) );
  INV_X4 U8112 ( .A(n6735), .ZN(n6738) );
  INV_X4 U8113 ( .A(n6735), .ZN(n6736) );
  INV_X4 U8114 ( .A(n6735), .ZN(n6737) );
  INV_X4 U8115 ( .A(n6739), .ZN(n6742) );
  INV_X4 U8116 ( .A(n6739), .ZN(n6740) );
  INV_X4 U8117 ( .A(n6739), .ZN(n6741) );
  INV_X4 U8118 ( .A(n6746), .ZN(n6747) );
  INV_X4 U8119 ( .A(n6746), .ZN(n6748) );
  INV_X4 U8120 ( .A(n340), .ZN(n6754) );
  INV_X4 U8121 ( .A(n6754), .ZN(n6753) );
  INV_X4 U8122 ( .A(n6754), .ZN(n6752) );
  INV_X4 U8123 ( .A(n5297), .ZN(n6755) );
  INV_X4 U8124 ( .A(n5297), .ZN(n6756) );
  INV_X4 U8125 ( .A(n5298), .ZN(n6758) );
  INV_X4 U8126 ( .A(n5298), .ZN(n6759) );
  INV_X4 U8127 ( .A(n5290), .ZN(n6769) );
  INV_X4 U8128 ( .A(n5290), .ZN(n6768) );
  INV_X4 U8129 ( .A(n6771), .ZN(n6774) );
  INV_X4 U8130 ( .A(n6771), .ZN(n6772) );
  INV_X4 U8131 ( .A(n6771), .ZN(n6773) );
  INV_X4 U8132 ( .A(n6692), .ZN(n6695) );
  INV_X4 U8133 ( .A(n6692), .ZN(n6693) );
  INV_X4 U8134 ( .A(n6692), .ZN(n6694) );
  INV_X4 U8135 ( .A(n5300), .ZN(n6689) );
  INV_X4 U8136 ( .A(n5300), .ZN(n6690) );
  INV_X2 U8137 ( .A(n5309), .ZN(n10101) );
  INV_X4 U8138 ( .A(n6696), .ZN(n6697) );
  INV_X4 U8139 ( .A(n6696), .ZN(n6698) );
  INV_X4 U8140 ( .A(n6696), .ZN(n6699) );
  INV_X16 U8141 ( .A(n6514), .ZN(n6515) );
  INV_X2 U8142 ( .A(n6515), .ZN(n11812) );
  INV_X2 U8143 ( .A(n6568), .ZN(n5916) );
  INV_X4 U8144 ( .A(net368201), .ZN(net375435) );
  NAND2_X2 U8145 ( .A1(n9188), .A2(n9189), .ZN(n13222) );
  OR2_X4 U8146 ( .A1(aluBoi_aluBoi_shft_sraout[21]), .A2(
        aluBoi_aluBoi_shft_sraout[20]), .ZN(n5717) );
  INV_X4 U8147 ( .A(regRst), .ZN(n6958) );
  INV_X4 U8148 ( .A(regRst), .ZN(n6957) );
  INV_X4 U8149 ( .A(regRst), .ZN(n6956) );
  INV_X4 U8150 ( .A(regRst), .ZN(n6955) );
  OR2_X4 U8151 ( .A1(n13199), .A2(n13151), .ZN(n5718) );
  OR2_X4 U8152 ( .A1(aluBoi_aluBoi_shft_sllout[19]), .A2(
        aluBoi_aluBoi_shft_sllout[18]), .ZN(n5719) );
  INV_X4 U8153 ( .A(pcRst), .ZN(n6961) );
  INV_X4 U8154 ( .A(pcRst), .ZN(n6960) );
  NAND2_X1 U8155 ( .A1(aluBoi_imm32w_4_), .A2(n6556), .ZN(n8230) );
  AOI222_X2 U8156 ( .A1(n13019), .A2(n13130), .B1(aluBoi_multBoi_temppp[17]), 
        .B2(net368069), .C1(n5316), .C2(aluBoi_imm32w_4_), .ZN(n13135) );
  XNOR2_X1 U8157 ( .A(n10360), .B(n10359), .ZN(n10362) );
  AOI22_X1 U8158 ( .A1(n6570), .A2(idOut_105_), .B1(n5751), .B2(n10165), .ZN(
        n5721) );
  XOR2_X1 U8159 ( .A(idOut_86_), .B(aluBoi_imm32w_0_), .Z(n10405) );
  NAND2_X1 U8160 ( .A1(aluBoi_imm32w_0_), .A2(n6556), .ZN(n8709) );
  AOI22_X1 U8161 ( .A1(n10126), .A2(n9928), .B1(ifOut_86_), .B2(ifInst[22]), 
        .ZN(n5722) );
  BUF_X32 U8162 ( .A(n10085), .Z(n5723) );
  XOR2_X2 U8163 ( .A(n5725), .B(n6073), .Z(n5724) );
  INV_X4 U8164 ( .A(n5724), .ZN(n10386) );
  BUF_X32 U8165 ( .A(n10295), .Z(n5726) );
  NAND2_X4 U8166 ( .A1(iaddr[21]), .A2(n10144), .ZN(n12710) );
  BUF_X32 U8167 ( .A(n10322), .Z(n5727) );
  XNOR2_X2 U8168 ( .A(n5728), .B(n6079), .ZN(n9203) );
  INV_X1 U8169 ( .A(n10291), .ZN(n5729) );
  INV_X4 U8170 ( .A(n5729), .ZN(n5730) );
  AOI22_X1 U8171 ( .A1(n10150), .A2(n9926), .B1(ifOut_84_), .B2(ifInst[20]), 
        .ZN(n5731) );
  INV_X1 U8172 ( .A(n13152), .ZN(n9204) );
  BUF_X32 U8173 ( .A(n10243), .Z(n5733) );
  OAI21_X2 U8174 ( .B1(n10035), .B2(n10332), .A(n6548), .ZN(n10036) );
  OAI21_X2 U8175 ( .B1(n10299), .B2(n10332), .A(n10298), .ZN(n10301) );
  NOR2_X1 U8176 ( .A1(iaddr[5]), .A2(n10332), .ZN(n10333) );
  BUF_X32 U8177 ( .A(n10351), .Z(n5734) );
  BUF_X32 U8178 ( .A(n10268), .Z(n5735) );
  AOI222_X2 U8179 ( .A1(n13019), .A2(n13112), .B1(aluBoi_multBoi_temppp[14]), 
        .B2(net368069), .C1(n5316), .C2(aluBoi_imm32w_1_), .ZN(n13117) );
  XNOR2_X1 U8180 ( .A(idOut_87_), .B(aluBoi_imm32w_1_), .ZN(n10394) );
  OAI21_X2 U8181 ( .B1(n13182), .B2(n13181), .A(n13062), .ZN(n13184) );
  AOI22_X1 U8182 ( .A1(n10228), .A2(n9920), .B1(ifOut_78_), .B2(ifInst[14]), 
        .ZN(n5736) );
  BUF_X32 U8183 ( .A(n10167), .Z(n5737) );
  NAND2_X2 U8184 ( .A1(n6571), .A2(n12687), .ZN(n10102) );
  NAND2_X4 U8185 ( .A1(n9986), .A2(iaddr[23]), .ZN(n12687) );
  OAI211_X4 U8186 ( .C1(n9203), .C2(n13222), .A(n9202), .B(n9201), .ZN(n13152)
         );
  AOI22_X1 U8187 ( .A1(n10210), .A2(n9922), .B1(ifOut_80_), .B2(ifInst[16]), 
        .ZN(n5738) );
  AOI22_X1 U8188 ( .A1(n10339), .A2(n9912), .B1(ifOut_70_), .B2(ifInst[6]), 
        .ZN(n5739) );
  AOI22_X1 U8189 ( .A1(n10278), .A2(n9916), .B1(ifOut_74_), .B2(ifInst[10]), 
        .ZN(n5740) );
  BUF_X32 U8190 ( .A(n5755), .Z(n5741) );
  INV_X2 U8191 ( .A(n13049), .ZN(n13050) );
  AOI22_X1 U8192 ( .A1(n10253), .A2(n9918), .B1(ifOut_76_), .B2(ifInst[12]), 
        .ZN(n5742) );
  XNOR2_X1 U8193 ( .A(n10378), .B(n10377), .ZN(n10379) );
  INV_X8 U8194 ( .A(n12805), .ZN(n10239) );
  AOI21_X1 U8195 ( .B1(n10286), .B2(n12805), .A(n6434), .ZN(n10240) );
  NAND2_X4 U8196 ( .A1(iaddr[12]), .A2(n10259), .ZN(n12805) );
  XNOR2_X1 U8197 ( .A(n5723), .B(n10084), .ZN(n10097) );
  INV_X4 U8198 ( .A(n10592), .ZN(n5743) );
  OAI22_X4 U8199 ( .A1(net362107), .A2(net362108), .B1(net362110), .B2(
        net362109), .ZN(n10592) );
  INV_X2 U8200 ( .A(n10592), .ZN(n10595) );
  XNOR2_X1 U8201 ( .A(n5731), .B(n10137), .ZN(n10140) );
  XNOR2_X1 U8202 ( .A(n5722), .B(n10112), .ZN(n10120) );
  INV_X1 U8203 ( .A(n5721), .ZN(n10152) );
  XNOR2_X1 U8204 ( .A(n10326), .B(n5739), .ZN(n10327) );
  XNOR2_X1 U8205 ( .A(n10272), .B(n5740), .ZN(n10273) );
  XNOR2_X1 U8206 ( .A(n10387), .B(n10386), .ZN(n10388) );
  XNOR2_X1 U8207 ( .A(n5733), .B(n10244), .ZN(n10249) );
  XNOR2_X1 U8208 ( .A(n10247), .B(n5742), .ZN(n10248) );
  XNOR2_X1 U8209 ( .A(n10222), .B(n5736), .ZN(n10223) );
  OAI22_X1 U8210 ( .A1(n6568), .A2(n5486), .B1(n10175), .B2(n5741), .ZN(n5746)
         );
  INV_X1 U8211 ( .A(n5741), .ZN(n10176) );
  XNOR2_X1 U8212 ( .A(n10385), .B(n10384), .ZN(n10389) );
  INV_X2 U8213 ( .A(n5915), .ZN(n10087) );
  INV_X1 U8214 ( .A(n9975), .ZN(n5744) );
  BUF_X16 U8215 ( .A(n5017), .Z(n5745) );
  INV_X8 U8216 ( .A(n10061), .ZN(n9975) );
  AOI21_X1 U8217 ( .B1(n10286), .B2(n12730), .A(n6434), .ZN(n10157) );
  NAND2_X4 U8218 ( .A1(iaddr[19]), .A2(n10161), .ZN(n12730) );
  INV_X1 U8219 ( .A(n9968), .ZN(n5747) );
  INV_X8 U8220 ( .A(n10128), .ZN(n9968) );
  OAI21_X4 U8221 ( .B1(n10291), .B2(n10292), .A(n9915), .ZN(n10278) );
  AOI22_X4 U8222 ( .A1(n10306), .A2(n9914), .B1(ifOut_72_), .B2(ifInst[8]), 
        .ZN(n10291) );
  BUF_X32 U8223 ( .A(n13210), .Z(n5748) );
  OAI21_X2 U8224 ( .B1(n13210), .B2(n13209), .A(n13062), .ZN(n13212) );
  OAI211_X4 U8225 ( .C1(n9739), .C2(n13222), .A(n9738), .B(n9737), .ZN(n13210)
         );
  INV_X8 U8226 ( .A(n12791), .ZN(n10234) );
  AOI21_X1 U8227 ( .B1(n10286), .B2(n12791), .A(n6434), .ZN(n10235) );
  NAND2_X4 U8228 ( .A1(iaddr[13]), .A2(n10239), .ZN(n12791) );
  OAI21_X4 U8229 ( .B1(n10167), .B2(n10166), .A(n9925), .ZN(n10150) );
  AOI22_X4 U8230 ( .A1(n10174), .A2(n9924), .B1(ifOut_82_), .B2(ifInst[18]), 
        .ZN(n10167) );
  NAND2_X1 U8231 ( .A1(n6590), .A2(aluBoi_imm32w_0_), .ZN(n13413) );
  AOI222_X2 U8232 ( .A1(n12982), .A2(n13123), .B1(aluBoi_multBoi_temppp[13]), 
        .B2(net368069), .C1(n5316), .C2(aluBoi_imm32w_0_), .ZN(n13128) );
  NAND2_X4 U8233 ( .A1(idOut_86_), .A2(aluBoi_imm32w_0_), .ZN(n10392) );
  BUF_X4 U8234 ( .A(n10374), .Z(n5754) );
  AOI22_X4 U8235 ( .A1(n10387), .A2(n5724), .B1(idOut_88_), .B2(
        aluBoi_imm32w_2_), .ZN(n10374) );
  OAI21_X4 U8236 ( .B1(n10193), .B2(n10192), .A(n9923), .ZN(n10174) );
  AOI22_X4 U8237 ( .A1(n10210), .A2(n9922), .B1(ifOut_80_), .B2(ifInst[16]), 
        .ZN(n10193) );
  INV_X1 U8238 ( .A(n12969), .ZN(n12972) );
  AOI22_X4 U8239 ( .A1(n6570), .A2(idOut_105_), .B1(n5751), .B2(n10165), .ZN(
        n5750) );
  INV_X4 U8240 ( .A(n6570), .ZN(n6569) );
  NAND2_X1 U8241 ( .A1(iaddr[3]), .A2(n6604), .ZN(n12891) );
  NAND2_X1 U8242 ( .A1(iaddr[3]), .A2(iaddr[2]), .ZN(n12883) );
  NAND2_X4 U8243 ( .A1(iaddr[4]), .A2(iaddr[3]), .ZN(n12876) );
  AOI21_X1 U8244 ( .B1(n10286), .B2(n12786), .A(n6434), .ZN(n10216) );
  INV_X1 U8245 ( .A(n12786), .ZN(n12771) );
  NAND2_X4 U8246 ( .A1(iaddr[14]), .A2(n10234), .ZN(n12786) );
  INV_X2 U8247 ( .A(n10373), .ZN(n10375) );
  OAI21_X2 U8248 ( .B1(n13200), .B2(n13199), .A(n13062), .ZN(n13202) );
  OAI221_X2 U8249 ( .B1(n9766), .B2(n9754), .C1(n9753), .C2(n13222), .A(n9752), 
        .ZN(n13200) );
  OAI21_X4 U8250 ( .B1(n10348), .B2(n10347), .A(n9911), .ZN(n10339) );
  AOI22_X4 U8251 ( .A1(n10358), .A2(n9910), .B1(ifOut_68_), .B2(ifInst[4]), 
        .ZN(n10348) );
  INV_X4 U8252 ( .A(n5912), .ZN(n10667) );
  NOR2_X4 U8253 ( .A1(net367631), .A2(n12326), .ZN(aluBoi_multBoi_N49) );
  NAND2_X2 U8254 ( .A1(net359554), .A2(net359555), .ZN(net359785) );
  NOR3_X1 U8255 ( .A1(n5748), .A2(n13238), .A3(n13200), .ZN(n9773) );
  AOI22_X4 U8256 ( .A1(n10100), .A2(n5352), .B1(ifOut_88_), .B2(ifInst[24]), 
        .ZN(n10085) );
  NAND2_X4 U8257 ( .A1(n12221), .A2(net359923), .ZN(n12324) );
  NAND2_X4 U8258 ( .A1(n10881), .A2(net361709), .ZN(n12221) );
  NOR2_X1 U8259 ( .A1(net359554), .A2(net359555), .ZN(net359552) );
  NAND2_X1 U8260 ( .A1(aluBoi_multBoi_temppp[36]), .A2(n6045), .ZN(n10872) );
  XOR2_X2 U8261 ( .A(n9380), .B(n9376), .Z(n9187) );
  AOI22_X4 U8262 ( .A1(n10126), .A2(n9928), .B1(ifOut_86_), .B2(ifInst[22]), 
        .ZN(n10113) );
  NAND2_X1 U8263 ( .A1(n9741), .A2(n9740), .ZN(n5753) );
  AOI22_X4 U8264 ( .A1(n5756), .A2(idOut_103_), .B1(n5757), .B2(n10191), .ZN(
        n5755) );
  INV_X4 U8265 ( .A(n9081), .ZN(n8882) );
  OAI21_X1 U8266 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9092) );
  INV_X8 U8267 ( .A(n5993), .ZN(n8706) );
  OAI22_X4 U8268 ( .A1(n13269), .A2(n6036), .B1(n5994), .B2(n5714), .ZN(n5993)
         );
  INV_X1 U8269 ( .A(n9103), .ZN(n9108) );
  OAI21_X1 U8270 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9079) );
  INV_X8 U8271 ( .A(n12640), .ZN(n10035) );
  NOR2_X1 U8272 ( .A1(n12640), .A2(n6551), .ZN(n10037) );
  OAI211_X1 U8273 ( .C1(iaddr[28]), .C2(n9987), .A(n12640), .B(n6603), .ZN(
        n12642) );
  NAND2_X4 U8274 ( .A1(iaddr[28]), .A2(n9987), .ZN(n12640) );
  INV_X8 U8275 ( .A(n12625), .ZN(n10010) );
  OAI211_X1 U8276 ( .C1(iaddr[29]), .C2(n10035), .A(n12625), .B(n6603), .ZN(
        n12627) );
  NAND2_X4 U8277 ( .A1(iaddr[29]), .A2(n10035), .ZN(n12625) );
  OAI211_X2 U8278 ( .C1(n9985), .C2(n9984), .A(n9983), .B(n6576), .ZN(n9998)
         );
  OAI211_X1 U8279 ( .C1(n5019), .C2(n13375), .A(n13268), .B(n13267), .ZN(
        n13659) );
  MUX2_X1 U8280 ( .A(n8348), .B(n8347), .S(n6808), .Z(n8349) );
  MUX2_X1 U8281 ( .A(n8352), .B(n8351), .S(n6831), .Z(n8353) );
  INV_X8 U8282 ( .A(net378138), .ZN(n5763) );
  MUX2_X2 U8283 ( .A(regBoiz_regfile_30__31_), .B(regBoiz_regfile_31__31_), 
        .S(net369156), .Z(n8347) );
  MUX2_X1 U8284 ( .A(n8350), .B(n8349), .S(n6826), .Z(n8351) );
  INV_X16 U8285 ( .A(n6615), .ZN(n6614) );
  NAND2_X1 U8286 ( .A1(idOut_88_), .A2(n6588), .ZN(n12900) );
  INV_X16 U8287 ( .A(net369158), .ZN(net369232) );
  INV_X32 U8288 ( .A(net378138), .ZN(net369160) );
  MUX2_X2 U8289 ( .A(n5759), .B(n5760), .S(net369240), .Z(n5758) );
  MUX2_X1 U8290 ( .A(n8320), .B(n8319), .S(n6826), .Z(n8321) );
  MUX2_X2 U8291 ( .A(n8309), .B(n8310), .S(n6815), .Z(n8314) );
  XNOR2_X1 U8292 ( .A(n10375), .B(n5754), .ZN(n10380) );
  XNOR2_X1 U8293 ( .A(n5747), .B(n10127), .ZN(n10129) );
  XNOR2_X2 U8294 ( .A(n10754), .B(net362026), .ZN(n5761) );
  INV_X4 U8295 ( .A(n10862), .ZN(n6056) );
  AOI22_X4 U8296 ( .A1(n10150), .A2(n9926), .B1(ifOut_84_), .B2(ifInst[20]), 
        .ZN(n10138) );
  NAND2_X2 U8297 ( .A1(n11917), .A2(n11953), .ZN(n11959) );
  NAND2_X2 U8298 ( .A1(n9745), .A2(n13220), .ZN(n9748) );
  INV_X8 U8299 ( .A(n13709), .ZN(n6615) );
  NAND2_X4 U8300 ( .A1(n5927), .A2(n13219), .ZN(n9727) );
  XNOR2_X2 U8301 ( .A(n8701), .B(n5762), .ZN(n5955) );
  INV_X2 U8302 ( .A(n8699), .ZN(n6038) );
  XNOR2_X1 U8303 ( .A(n10323), .B(n5727), .ZN(n10328) );
  AOI22_X4 U8304 ( .A1(n10337), .A2(n9953), .B1(idOut_92_), .B2(
        aluBoi_imm32w_6_), .ZN(n10322) );
  AOI22_X4 U8305 ( .A1(n10280), .A2(n9957), .B1(idOut_96_), .B2(
        aluBoi_imm32w_10_), .ZN(n10268) );
  AOI211_X2 U8306 ( .C1(n5753), .C2(n9761), .A(n9744), .B(n9743), .ZN(n9749)
         );
  NAND2_X4 U8307 ( .A1(n10010), .A2(iaddr[30]), .ZN(n12613) );
  XNOR2_X1 U8308 ( .A(n5744), .B(n10060), .ZN(n10062) );
  XNOR2_X1 U8309 ( .A(n10269), .B(n5735), .ZN(n10274) );
  AOI22_X4 U8310 ( .A1(n10228), .A2(n9920), .B1(ifOut_78_), .B2(ifInst[14]), 
        .ZN(n10221) );
  XNOR2_X1 U8311 ( .A(n10352), .B(n5734), .ZN(n10353) );
  AOI22_X4 U8312 ( .A1(n10360), .A2(n9951), .B1(idOut_90_), .B2(
        aluBoi_imm32w_4_), .ZN(n10351) );
  XOR2_X1 U8313 ( .A(n10296), .B(n5726), .Z(n10297) );
  AOI22_X4 U8314 ( .A1(n10308), .A2(n9955), .B1(idOut_94_), .B2(
        aluBoi_imm32w_8_), .ZN(n10295) );
  NOR3_X1 U8315 ( .A1(n13182), .A2(n13192), .A3(n13172), .ZN(n9772) );
  OAI221_X4 U8316 ( .B1(n9766), .B2(n9765), .C1(n9764), .C2(n13222), .A(n9763), 
        .ZN(n13192) );
  OAI21_X2 U8317 ( .B1(n13194), .B2(n13231), .A(n13193), .ZN(n4765) );
  OAI21_X4 U8318 ( .B1(n12249), .B2(n9456), .A(n9745), .ZN(n5927) );
  NAND3_X2 U8319 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n13709) );
  NAND2_X2 U8320 ( .A1(n9085), .A2(n9086), .ZN(n8714) );
  AOI22_X4 U8321 ( .A1(n10278), .A2(n9916), .B1(ifOut_74_), .B2(ifInst[10]), 
        .ZN(n10271) );
  XNOR2_X1 U8322 ( .A(n10176), .B(n10175), .ZN(n10179) );
  XNOR2_X1 U8323 ( .A(n5746), .B(n10164), .ZN(n10170) );
  INV_X4 U8324 ( .A(net369232), .ZN(net369230) );
  INV_X4 U8325 ( .A(n8699), .ZN(n6037) );
  NAND2_X1 U8326 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  NAND3_X2 U8327 ( .A1(n8661), .A2(n8660), .A3(n8659), .ZN(n10416) );
  INV_X16 U8328 ( .A(net369232), .ZN(net369228) );
  INV_X16 U8329 ( .A(net369232), .ZN(net369226) );
  NAND3_X2 U8330 ( .A1(n8695), .A2(n8694), .A3(n8693), .ZN(n10412) );
  NAND2_X1 U8331 ( .A1(n8930), .A2(n8883), .ZN(n8766) );
  MUX2_X1 U8332 ( .A(regBoiz_regfile_30__26_), .B(regBoiz_regfile_31__26_), 
        .S(net369165), .Z(n8685) );
  MUX2_X1 U8333 ( .A(regBoiz_regfile_14__23_), .B(regBoiz_regfile_15__23_), 
        .S(net369165), .Z(n8527) );
  MUX2_X2 U8334 ( .A(regBoiz_regfile_14__22_), .B(regBoiz_regfile_15__22_), 
        .S(net369161), .Z(n8597) );
  MUX2_X1 U8335 ( .A(regBoiz_regfile_10__22_), .B(regBoiz_regfile_11__22_), 
        .S(net369166), .Z(n8595) );
  INV_X32 U8336 ( .A(net369160), .ZN(net369165) );
  NAND2_X2 U8337 ( .A1(n9718), .A2(n13036), .ZN(n8660) );
  INV_X1 U8338 ( .A(n13036), .ZN(n13039) );
  OAI211_X2 U8339 ( .C1(n12506), .C2(n12505), .A(n5025), .B(net100619), .ZN(
        n12507) );
  OAI22_X4 U8340 ( .A1(n6568), .A2(n5486), .B1(n5755), .B2(n10175), .ZN(n10165) );
  NOR3_X1 U8341 ( .A1(n5462), .A2(idOut_115_), .A3(n5017), .ZN(n10032) );
  XNOR2_X1 U8342 ( .A(n5745), .B(n10044), .ZN(n10056) );
  AOI22_X4 U8343 ( .A1(n10339), .A2(n9912), .B1(ifOut_70_), .B2(ifInst[6]), 
        .ZN(n10325) );
  OAI211_X1 U8344 ( .C1(net361260), .C2(net361261), .A(n11364), .B(net100619), 
        .ZN(n11170) );
  INV_X4 U8345 ( .A(net359915), .ZN(net360914) );
  NOR2_X2 U8346 ( .A1(net359553), .A2(net359784), .ZN(net359782) );
  XNOR2_X2 U8347 ( .A(net359782), .B(n5223), .ZN(n12326) );
  NAND2_X4 U8348 ( .A1(net359550), .A2(n12502), .ZN(n12501) );
  INV_X4 U8349 ( .A(n11951), .ZN(n6013) );
  NOR3_X2 U8350 ( .A1(n5418), .A2(n11952), .A3(n11951), .ZN(n11950) );
  INV_X8 U8351 ( .A(n11947), .ZN(n11951) );
  AOI21_X2 U8352 ( .B1(n11370), .B2(n12328), .A(net360915), .ZN(n11438) );
  AOI22_X4 U8353 ( .A1(n10253), .A2(n9918), .B1(ifOut_76_), .B2(ifInst[12]), 
        .ZN(n10246) );
  NOR2_X2 U8354 ( .A1(n12231), .A2(net367631), .ZN(aluBoi_multBoi_N63) );
  XNOR2_X1 U8355 ( .A(n10152), .B(n10151), .ZN(n10154) );
  INV_X4 U8356 ( .A(n10099), .ZN(n5917) );
  NAND2_X2 U8357 ( .A1(n5767), .A2(n12982), .ZN(n13515) );
  NOR3_X2 U8358 ( .A1(n13222), .A2(n13221), .A3(n5927), .ZN(n13229) );
  XOR2_X1 U8359 ( .A(n10292), .B(n5730), .Z(n10294) );
  NAND3_X4 U8360 ( .A1(net377817), .A2(net377791), .A3(
        aluBoi_multBoi_temppp[49]), .ZN(net359533) );
  OAI21_X2 U8361 ( .B1(n6625), .B2(n6726), .A(n654), .ZN(n4412) );
  AOI21_X4 U8362 ( .B1(n12229), .B2(n12519), .A(n12228), .ZN(n12230) );
  INV_X1 U8363 ( .A(n9780), .ZN(n5765) );
  INV_X4 U8364 ( .A(n5765), .ZN(n5766) );
  XNOR2_X2 U8365 ( .A(n9780), .B(n5768), .ZN(n5767) );
  OAI21_X2 U8366 ( .B1(n9082), .B2(n5018), .A(n9080), .ZN(n9084) );
  XNOR2_X2 U8367 ( .A(n8702), .B(n8701), .ZN(n9081) );
  INV_X16 U8368 ( .A(net369158), .ZN(net369216) );
  INV_X32 U8369 ( .A(net369139), .ZN(net369144) );
  NOR2_X1 U8370 ( .A1(net359680), .A2(n11971), .ZN(n11973) );
  BUF_X4 U8371 ( .A(net369138), .Z(net369142) );
  CLKBUF_X2 U8372 ( .A(n9105), .Z(n6052) );
  CLKBUF_X3 U8373 ( .A(n9116), .Z(n5978) );
  NAND2_X2 U8374 ( .A1(n12225), .A2(n12509), .ZN(n12226) );
  NAND2_X1 U8375 ( .A1(n10994), .A2(n10999), .ZN(n11102) );
  OAI21_X2 U8376 ( .B1(n10934), .B2(n10933), .A(n10999), .ZN(n10976) );
  OAI21_X2 U8377 ( .B1(n5657), .B2(n6734), .A(n596), .ZN(n4084) );
  INV_X8 U8378 ( .A(net361833), .ZN(net361832) );
  NAND2_X4 U8379 ( .A1(net361911), .A2(n10748), .ZN(net361833) );
  NAND2_X4 U8380 ( .A1(regBoiz_regfile_26__25_), .A2(n6787), .ZN(n7888) );
  OAI21_X2 U8381 ( .B1(n7891), .B2(n7890), .A(net366969), .ZN(n7892) );
  AOI21_X2 U8382 ( .B1(n7887), .B2(n7886), .A(net366951), .ZN(n7891) );
  AOI21_X2 U8383 ( .B1(n7889), .B2(n7888), .A(net366927), .ZN(n7890) );
  NAND3_X2 U8384 ( .A1(n11565), .A2(n11563), .A3(n11564), .ZN(n5772) );
  OAI21_X2 U8385 ( .B1(net377979), .B2(n12532), .A(n12339), .ZN(n12340) );
  NAND2_X4 U8386 ( .A1(n5773), .A2(net361387), .ZN(net361433) );
  INV_X8 U8387 ( .A(net361526), .ZN(net361387) );
  NAND2_X4 U8388 ( .A1(net361387), .A2(n5773), .ZN(net376785) );
  NAND3_X2 U8389 ( .A1(net361387), .A2(net369287), .A3(n5773), .ZN(net361386)
         );
  NAND2_X4 U8390 ( .A1(net375305), .A2(net361529), .ZN(net361526) );
  NAND3_X4 U8391 ( .A1(net361530), .A2(net361532), .A3(net377383), .ZN(
        net361529) );
  NOR2_X4 U8392 ( .A1(n5776), .A2(n5777), .ZN(net361530) );
  NAND2_X1 U8393 ( .A1(net378405), .A2(net361903), .ZN(n5778) );
  INV_X4 U8394 ( .A(net375304), .ZN(net375305) );
  NAND2_X2 U8395 ( .A1(n5782), .A2(net361539), .ZN(n5775) );
  INV_X4 U8396 ( .A(net361886), .ZN(net361539) );
  NOR2_X2 U8397 ( .A1(net361539), .A2(net361827), .ZN(net361825) );
  NAND4_X4 U8398 ( .A1(net361356), .A2(net376121), .A3(net361358), .A4(n5782), 
        .ZN(net361814) );
  NAND2_X1 U8399 ( .A1(net361358), .A2(n5782), .ZN(net361354) );
  INV_X8 U8400 ( .A(n5782), .ZN(net376691) );
  XNOR2_X2 U8401 ( .A(net361902), .B(net361537), .ZN(n5781) );
  NAND3_X2 U8402 ( .A1(net361524), .A2(net361437), .A3(net361523), .ZN(n5774)
         );
  NOR2_X4 U8403 ( .A1(net361541), .A2(n5779), .ZN(n5773) );
  XNOR2_X2 U8404 ( .A(net361543), .B(n5780), .ZN(n5779) );
  NAND2_X1 U8405 ( .A1(n5783), .A2(net361546), .ZN(n5780) );
  XNOR2_X2 U8406 ( .A(n10794), .B(n5783), .ZN(net361749) );
  INV_X8 U8407 ( .A(net361545), .ZN(net361629) );
  NAND3_X4 U8408 ( .A1(n5784), .A2(net376582), .A3(net360621), .ZN(net360609)
         );
  NAND3_X4 U8409 ( .A1(net360608), .A2(net360609), .A3(net359913), .ZN(
        net360284) );
  NOR3_X4 U8410 ( .A1(net360623), .A2(net360625), .A3(n5785), .ZN(n5784) );
  INV_X8 U8411 ( .A(n5789), .ZN(n5785) );
  NOR3_X2 U8412 ( .A1(n5785), .A2(net360634), .A3(net360635), .ZN(net360633)
         );
  NAND2_X4 U8413 ( .A1(aluBoi_multBoi_temppp[47]), .A2(n5790), .ZN(n5789) );
  INV_X4 U8414 ( .A(net360919), .ZN(n5790) );
  NAND2_X2 U8415 ( .A1(aluBoi_multBoi_temppp[47]), .A2(n5790), .ZN(net360996)
         );
  INV_X8 U8416 ( .A(net360626), .ZN(net360625) );
  NAND2_X4 U8417 ( .A1(n5786), .A2(net360628), .ZN(net360623) );
  NOR2_X4 U8418 ( .A1(net360629), .A2(n5787), .ZN(n5786) );
  INV_X4 U8419 ( .A(net360632), .ZN(net360629) );
  INV_X4 U8420 ( .A(net376581), .ZN(net376582) );
  NAND2_X1 U8421 ( .A1(net359915), .A2(net376582), .ZN(net359914) );
  NAND2_X4 U8422 ( .A1(aluBoi_multBoi_temppp[45]), .A2(n5791), .ZN(net360621)
         );
  NAND3_X2 U8423 ( .A1(net360633), .A2(net359916), .A3(net360621), .ZN(
        net360608) );
  OAI21_X4 U8424 ( .B1(net359918), .B2(net359919), .A(net360621), .ZN(
        net359550) );
  INV_X4 U8425 ( .A(n5788), .ZN(n5791) );
  INV_X8 U8426 ( .A(net361006), .ZN(net361000) );
  OAI21_X2 U8427 ( .B1(net361000), .B2(net361001), .A(net361002), .ZN(
        net378491) );
  NAND2_X4 U8428 ( .A1(net361007), .A2(net361008), .ZN(net361006) );
  NAND2_X2 U8429 ( .A1(net361025), .A2(n5793), .ZN(n5792) );
  INV_X4 U8430 ( .A(net361019), .ZN(n5793) );
  NAND2_X2 U8431 ( .A1(net360636), .A2(net360631), .ZN(net360635) );
  INV_X8 U8432 ( .A(net360628), .ZN(net360634) );
  NOR2_X2 U8433 ( .A1(net360915), .A2(net360634), .ZN(net360639) );
  NAND2_X2 U8434 ( .A1(net360605), .A2(net360604), .ZN(n5794) );
  NAND2_X4 U8435 ( .A1(net360007), .A2(net360008), .ZN(net360006) );
  NAND2_X4 U8436 ( .A1(net360005), .A2(net360006), .ZN(net359471) );
  NAND2_X4 U8437 ( .A1(n5804), .A2(n5795), .ZN(net360288) );
  INV_X8 U8438 ( .A(net360266), .ZN(n5795) );
  INV_X1 U8439 ( .A(n5795), .ZN(net378220) );
  NAND2_X2 U8440 ( .A1(n5022), .A2(n5795), .ZN(net359537) );
  INV_X4 U8441 ( .A(n5804), .ZN(net377342) );
  NOR3_X4 U8442 ( .A1(net359911), .A2(n5796), .A3(n5805), .ZN(net360287) );
  NAND2_X2 U8443 ( .A1(net359533), .A2(net359535), .ZN(n5805) );
  INV_X4 U8444 ( .A(net360273), .ZN(n5796) );
  XNOR2_X1 U8445 ( .A(net359911), .B(n5483), .ZN(net360583) );
  OAI21_X4 U8446 ( .B1(n5797), .B2(n5798), .A(n5799), .ZN(net360008) );
  NAND3_X2 U8447 ( .A1(n5800), .A2(net359532), .A3(net375993), .ZN(n5799) );
  NOR2_X4 U8448 ( .A1(net377342), .A2(net360266), .ZN(n5800) );
  OAI21_X2 U8449 ( .B1(n5801), .B2(n5802), .A(n5803), .ZN(n5798) );
  NAND2_X2 U8450 ( .A1(n5521), .A2(net360259), .ZN(n5803) );
  NAND2_X1 U8451 ( .A1(net360261), .A2(net360273), .ZN(n5802) );
  INV_X4 U8452 ( .A(net360262), .ZN(n5801) );
  NAND3_X4 U8453 ( .A1(n5145), .A2(net376826), .A3(n5806), .ZN(net361532) );
  INV_X1 U8454 ( .A(net378420), .ZN(net378060) );
  NOR3_X2 U8455 ( .A1(n5123), .A2(net361830), .A3(net361832), .ZN(net361829)
         );
  NAND2_X4 U8456 ( .A1(net362127), .A2(net376139), .ZN(net362092) );
  NAND3_X1 U8457 ( .A1(net362125), .A2(net376139), .A3(net362127), .ZN(
        net362091) );
  INV_X8 U8458 ( .A(net361834), .ZN(net361831) );
  XNOR2_X2 U8459 ( .A(net361906), .B(net361907), .ZN(net377383) );
  XNOR2_X2 U8460 ( .A(net377383), .B(net361893), .ZN(net362026) );
  XNOR2_X2 U8461 ( .A(net361900), .B(n5807), .ZN(net361535) );
  INV_X2 U8462 ( .A(net361535), .ZN(net361899) );
  INV_X4 U8463 ( .A(n5808), .ZN(n5807) );
  XNOR2_X2 U8464 ( .A(net361900), .B(n5807), .ZN(net361891) );
  XNOR2_X2 U8465 ( .A(net361949), .B(net362166), .ZN(n5808) );
  INV_X4 U8466 ( .A(net361536), .ZN(net362166) );
  INV_X4 U8467 ( .A(net362194), .ZN(net361900) );
  MUX2_X2 U8468 ( .A(net365091), .B(n5809), .S(net366973), .Z(net365090) );
  INV_X32 U8469 ( .A(net368770), .ZN(net366901) );
  INV_X16 U8470 ( .A(net368787), .ZN(net368770) );
  NAND2_X1 U8471 ( .A1(net366899), .A2(net366953), .ZN(net365284) );
  MUX2_X2 U8472 ( .A(net375769), .B(net368927), .S(net368770), .Z(net366184)
         );
  MUX2_X2 U8473 ( .A(regBoiz_regfile_2__27_), .B(regBoiz_regfile_3__27_), .S(
        net369164), .Z(net364764) );
  MUX2_X2 U8474 ( .A(regBoiz_regfile_10__27_), .B(regBoiz_regfile_11__27_), 
        .S(net369166), .Z(net364779) );
  OAI21_X4 U8475 ( .B1(net368185), .B2(net362028), .A(n5811), .ZN(net361536)
         );
  INV_X16 U8476 ( .A(n5812), .ZN(net377611) );
  INV_X8 U8477 ( .A(n5810), .ZN(n5812) );
  NAND2_X4 U8478 ( .A1(net362179), .A2(net362265), .ZN(n5810) );
  OAI22_X1 U8479 ( .A1(net360360), .A2(net368446), .B1(n4987), .B2(net368187), 
        .ZN(net360474) );
  INV_X8 U8480 ( .A(net368439), .ZN(net368440) );
  INV_X8 U8481 ( .A(net368440), .ZN(net368442) );
  INV_X8 U8482 ( .A(net368440), .ZN(net368444) );
  NAND2_X4 U8483 ( .A1(aluBoi_multOut[1]), .A2(n5304), .ZN(net368439) );
  NAND2_X4 U8484 ( .A1(net361416), .A2(net369287), .ZN(n5813) );
  INV_X4 U8485 ( .A(n5122), .ZN(net361400) );
  INV_X8 U8486 ( .A(net369285), .ZN(net369287) );
  INV_X8 U8487 ( .A(net361380), .ZN(net369285) );
  INV_X8 U8488 ( .A(net369285), .ZN(net369286) );
  NAND2_X4 U8489 ( .A1(net361630), .A2(net378336), .ZN(net361380) );
  INV_X1 U8490 ( .A(net361510), .ZN(net378336) );
  INV_X4 U8491 ( .A(net361511), .ZN(net361510) );
  XNOR2_X2 U8492 ( .A(net361509), .B(net361510), .ZN(net361443) );
  OAI22_X2 U8493 ( .A1(net361631), .A2(net368446), .B1(net368185), .B2(
        net361417), .ZN(net361511) );
  NAND2_X2 U8494 ( .A1(aluBoi_multOut[2]), .A2(n5319), .ZN(net359750) );
  OAI22_X2 U8495 ( .A1(net360205), .A2(net368442), .B1(net368187), .B2(
        net360206), .ZN(net360198) );
  OAI22_X2 U8496 ( .A1(net360723), .A2(net368442), .B1(net368187), .B2(
        net360403), .ZN(net360513) );
  NAND2_X4 U8497 ( .A1(net365090), .A2(net365089), .ZN(net365088) );
  NAND2_X2 U8498 ( .A1(net365087), .A2(net365088), .ZN(net362286) );
  NAND2_X4 U8499 ( .A1(net365087), .A2(net365088), .ZN(net377937) );
  INV_X4 U8500 ( .A(net363057), .ZN(net365089) );
  NAND2_X2 U8501 ( .A1(net365100), .A2(net365089), .ZN(net365099) );
  INV_X16 U8502 ( .A(net366993), .ZN(net366973) );
  INV_X8 U8503 ( .A(net366985), .ZN(net366993) );
  INV_X16 U8504 ( .A(net366993), .ZN(net366971) );
  MUX2_X2 U8505 ( .A(net364971), .B(net364970), .S(net366993), .Z(net362387)
         );
  INV_X32 U8506 ( .A(net366989), .ZN(net366985) );
  INV_X32 U8507 ( .A(net367011), .ZN(net366989) );
  INV_X16 U8508 ( .A(net366989), .ZN(net366987) );
  INV_X16 U8509 ( .A(net367013), .ZN(net367011) );
  INV_X16 U8510 ( .A(net368775), .ZN(net367013) );
  INV_X8 U8511 ( .A(net367013), .ZN(net367009) );
  INV_X4 U8512 ( .A(net368676), .ZN(net368775) );
  MUX2_X2 U8513 ( .A(regBoiz_regfile_0__27_), .B(regBoiz_regfile_8__27_), .S(
        net376330), .Z(net365091) );
  INV_X8 U8514 ( .A(net369210), .ZN(net376330) );
  INV_X4 U8515 ( .A(net362286), .ZN(net362268) );
  NAND2_X4 U8516 ( .A1(n5814), .A2(net365093), .ZN(net365087) );
  MUX2_X2 U8517 ( .A(net365095), .B(n5815), .S(net366973), .Z(n5814) );
  MUX2_X2 U8518 ( .A(regBoiz_regfile_6__27_), .B(regBoiz_regfile_14__27_), .S(
        net377109), .Z(n5815) );
  INV_X4 U8519 ( .A(net366907), .ZN(net377109) );
  INV_X8 U8520 ( .A(net366911), .ZN(net366907) );
  INV_X32 U8521 ( .A(net366911), .ZN(net366905) );
  MUX2_X2 U8522 ( .A(regBoiz_regfile_4__27_), .B(regBoiz_regfile_12__27_), .S(
        net376331), .Z(net365095) );
  INV_X16 U8523 ( .A(net369210), .ZN(net376331) );
  INV_X16 U8524 ( .A(net368903), .ZN(net369210) );
  INV_X16 U8525 ( .A(net368787), .ZN(net368903) );
  XNOR2_X2 U8526 ( .A(n5028), .B(aluBoi_multBoi_temppp[54]), .ZN(net375910) );
  INV_X1 U8527 ( .A(net359652), .ZN(net377602) );
  INV_X4 U8528 ( .A(net359490), .ZN(net359652) );
  AOI22_X4 U8529 ( .A1(net359492), .A2(net377784), .B1(net377784), .B2(
        net359493), .ZN(net359489) );
  NAND2_X2 U8530 ( .A1(net359494), .A2(net359495), .ZN(net359493) );
  INV_X4 U8531 ( .A(net359756), .ZN(net359494) );
  NAND2_X2 U8532 ( .A1(net359494), .A2(net359471), .ZN(net359574) );
  INV_X4 U8533 ( .A(n5817), .ZN(n5816) );
  NAND3_X2 U8534 ( .A1(net359499), .A2(net377452), .A3(net359495), .ZN(n5817)
         );
  XNOR2_X2 U8535 ( .A(n5818), .B(net359418), .ZN(net359490) );
  NAND2_X1 U8536 ( .A1(net359490), .A2(net359470), .ZN(net359577) );
  INV_X4 U8537 ( .A(net129670), .ZN(net359418) );
  NAND2_X4 U8538 ( .A1(net359449), .A2(net359450), .ZN(n5818) );
  OAI21_X4 U8539 ( .B1(net360003), .B2(net360004), .A(net359471), .ZN(
        net359492) );
  NAND2_X4 U8540 ( .A1(net359492), .A2(net359501), .ZN(net360002) );
  OAI21_X2 U8541 ( .B1(net368209), .B2(net362238), .A(net362237), .ZN(
        net362262) );
  INV_X32 U8542 ( .A(net368467), .ZN(net360821) );
  NAND2_X4 U8543 ( .A1(aluBoi_multBoi_runProd_0_), .A2(n5307), .ZN(net359966)
         );
  NAND2_X2 U8544 ( .A1(aluBoi_multOut[1]), .A2(n5307), .ZN(net359877) );
  NAND2_X1 U8545 ( .A1(net362265), .A2(net368548), .ZN(net362264) );
  INV_X16 U8546 ( .A(net368547), .ZN(net368548) );
  INV_X8 U8547 ( .A(net362266), .ZN(net368547) );
  NAND2_X2 U8548 ( .A1(net364904), .A2(n5821), .ZN(net362266) );
  INV_X4 U8549 ( .A(net364803), .ZN(n5820) );
  NOR2_X2 U8550 ( .A1(n5820), .A2(net364906), .ZN(net364905) );
  OAI21_X1 U8551 ( .B1(net362342), .B2(n5820), .A(net362253), .ZN(net362341)
         );
  NAND2_X4 U8552 ( .A1(net377481), .A2(net362268), .ZN(net362270) );
  NAND2_X4 U8553 ( .A1(daddr[4]), .A2(net362342), .ZN(net362265) );
  INV_X8 U8554 ( .A(net364941), .ZN(net362342) );
  NAND2_X4 U8555 ( .A1(net365335), .A2(net365336), .ZN(net364904) );
  NAND4_X2 U8556 ( .A1(net359472), .A2(net359471), .A3(net359470), .A4(
        net359473), .ZN(net359469) );
  NOR3_X4 U8557 ( .A1(n5272), .A2(net377071), .A3(n5822), .ZN(net360005) );
  NAND3_X2 U8558 ( .A1(net359767), .A2(net359905), .A3(net360011), .ZN(n5822)
         );
  INV_X2 U8559 ( .A(n5272), .ZN(net376321) );
  AOI21_X4 U8560 ( .B1(net361273), .B2(net361272), .A(net361274), .ZN(n5823)
         );
  INV_X4 U8561 ( .A(net361279), .ZN(net361274) );
  INV_X1 U8562 ( .A(net361274), .ZN(net377502) );
  NAND2_X2 U8563 ( .A1(net361275), .A2(net361276), .ZN(net361273) );
  NAND2_X4 U8564 ( .A1(net361273), .A2(net361272), .ZN(net361278) );
  NAND2_X4 U8565 ( .A1(net377550), .A2(net361057), .ZN(net361272) );
  NAND3_X4 U8566 ( .A1(net361320), .A2(net361272), .A3(net361053), .ZN(
        net361324) );
  XNOR2_X2 U8567 ( .A(net361081), .B(net361080), .ZN(net361279) );
  XNOR2_X1 U8568 ( .A(net361279), .B(aluBoi_multBoi_temppp[42]), .ZN(net361277) );
  NAND2_X4 U8569 ( .A1(net361275), .A2(net361276), .ZN(net361320) );
  NAND2_X2 U8570 ( .A1(net361057), .A2(net361056), .ZN(net361088) );
  AND2_X2 U8571 ( .A1(net361056), .A2(net361057), .ZN(net375793) );
  INV_X4 U8572 ( .A(net361057), .ZN(net361342) );
  INV_X2 U8573 ( .A(net361081), .ZN(net361079) );
  NAND2_X2 U8574 ( .A1(net361409), .A2(net361081), .ZN(net361322) );
  NOR2_X2 U8575 ( .A1(net361079), .A2(net361080), .ZN(net361077) );
  NAND3_X4 U8576 ( .A1(net361411), .A2(net361410), .A3(net361080), .ZN(
        net361053) );
  INV_X4 U8577 ( .A(net361080), .ZN(net361409) );
  OAI211_X2 U8578 ( .C1(net359492), .C2(n5101), .A(net359462), .B(net359682), 
        .ZN(net359809) );
  NOR3_X4 U8579 ( .A1(net360015), .A2(n5825), .A3(n5824), .ZN(net360004) );
  XNOR2_X2 U8580 ( .A(net359899), .B(n5348), .ZN(n5824) );
  NAND2_X4 U8581 ( .A1(net360033), .A2(n5348), .ZN(net376916) );
  XNOR2_X2 U8582 ( .A(net359899), .B(n5348), .ZN(net359765) );
  NOR2_X4 U8583 ( .A1(net360014), .A2(net359504), .ZN(n5825) );
  NOR3_X4 U8584 ( .A1(n5827), .A2(net362114), .A3(n5834), .ZN(n5828) );
  OAI21_X4 U8585 ( .B1(n5828), .B2(n5829), .A(net377530), .ZN(net361834) );
  INV_X8 U8586 ( .A(n5833), .ZN(n5834) );
  NOR2_X4 U8587 ( .A1(n5827), .A2(n5834), .ZN(net362107) );
  INV_X8 U8588 ( .A(net362116), .ZN(n5833) );
  XNOR2_X2 U8589 ( .A(n5827), .B(n5833), .ZN(net362016) );
  NOR2_X2 U8590 ( .A1(net362114), .A2(net378432), .ZN(n5829) );
  NAND2_X2 U8591 ( .A1(net378432), .A2(net362114), .ZN(net362108) );
  XNOR2_X2 U8592 ( .A(net362321), .B(net362130), .ZN(n5826) );
  NAND2_X4 U8593 ( .A1(net362312), .A2(net362311), .ZN(net362116) );
  NAND2_X2 U8594 ( .A1(net362113), .A2(net362116), .ZN(net362121) );
  XNOR2_X2 U8595 ( .A(net362135), .B(net362136), .ZN(net362120) );
  NAND2_X2 U8596 ( .A1(net362121), .A2(net362120), .ZN(net362110) );
  NAND2_X4 U8597 ( .A1(n5832), .A2(net362051), .ZN(net362136) );
  NAND3_X2 U8598 ( .A1(net362139), .A2(net362063), .A3(net362138), .ZN(n5832)
         );
  XNOR2_X2 U8599 ( .A(net362231), .B(net362232), .ZN(net378103) );
  NAND2_X4 U8600 ( .A1(net362131), .A2(net362323), .ZN(net362321) );
  XNOR2_X2 U8601 ( .A(net362321), .B(net362130), .ZN(net377355) );
  NAND3_X2 U8602 ( .A1(n5831), .A2(net362052), .A3(net362049), .ZN(net362323)
         );
  INV_X8 U8603 ( .A(net362134), .ZN(n5831) );
  AOI21_X4 U8604 ( .B1(net362061), .B2(n5831), .A(net362196), .ZN(net362161)
         );
  AOI21_X4 U8605 ( .B1(net362061), .B2(n5831), .A(net362196), .ZN(net375794)
         );
  NAND3_X1 U8606 ( .A1(net362049), .A2(n5831), .A3(net362052), .ZN(n5830) );
  OAI22_X1 U8607 ( .A1(net362322), .A2(net359986), .B1(net362105), .B2(
        net368187), .ZN(net362130) );
  NAND3_X2 U8608 ( .A1(net362130), .A2(net362131), .A3(n5830), .ZN(net362113)
         );
  AOI21_X4 U8609 ( .B1(net361265), .B2(net361266), .A(net359783), .ZN(
        net361264) );
  OAI21_X4 U8610 ( .B1(net361263), .B2(net361262), .A(net361264), .ZN(
        net360626) );
  INV_X4 U8611 ( .A(net359554), .ZN(net361265) );
  XNOR2_X2 U8612 ( .A(net361268), .B(n5685), .ZN(net359783) );
  NAND3_X4 U8613 ( .A1(net361324), .A2(net361322), .A3(n5836), .ZN(net361271)
         );
  NAND3_X1 U8614 ( .A1(net361322), .A2(n5836), .A3(n5225), .ZN(net377660) );
  NOR2_X4 U8615 ( .A1(n5835), .A2(n5596), .ZN(net359784) );
  XNOR2_X2 U8616 ( .A(net377502), .B(net361278), .ZN(n5835) );
  XNOR2_X2 U8617 ( .A(net361277), .B(net361278), .ZN(net359554) );
  NAND3_X1 U8618 ( .A1(aluBoi_multBoi_temppp[43]), .A2(net361321), .A3(
        net377660), .ZN(net360632) );
  INV_X4 U8619 ( .A(net361270), .ZN(net361327) );
  NAND4_X4 U8620 ( .A1(net361322), .A2(net361319), .A3(net361318), .A4(
        net361335), .ZN(net361015) );
  NAND2_X2 U8621 ( .A1(net361322), .A2(n5836), .ZN(net361361) );
  NAND2_X4 U8622 ( .A1(net362146), .A2(net362140), .ZN(net361913) );
  NAND2_X2 U8623 ( .A1(aluBoi_multBoi_temppp[0]), .A2(n5304), .ZN(net359601)
         );
  OAI22_X2 U8624 ( .A1(n10570), .A2(net368436), .B1(net368181), .B2(net362124), 
        .ZN(net362096) );
  INV_X16 U8625 ( .A(net368501), .ZN(net376602) );
  INV_X8 U8626 ( .A(net334218), .ZN(net368501) );
  NAND2_X2 U8627 ( .A1(net377375), .A2(net361053), .ZN(net361270) );
  XNOR2_X2 U8628 ( .A(n5837), .B(net361394), .ZN(net361325) );
  INV_X4 U8629 ( .A(n5838), .ZN(n5837) );
  XNOR2_X2 U8630 ( .A(n5837), .B(net361394), .ZN(net377375) );
  XNOR2_X2 U8631 ( .A(n5837), .B(net361083), .ZN(net361076) );
  XNOR2_X2 U8632 ( .A(net361391), .B(net361372), .ZN(n5838) );
  INV_X4 U8633 ( .A(net377373), .ZN(net361372) );
  INV_X4 U8634 ( .A(net377375), .ZN(net361335) );
  OAI221_X4 U8635 ( .B1(net368215), .B2(net362233), .C1(n5840), .C2(n5841), 
        .A(n5842), .ZN(net362232) );
  XOR2_X2 U8636 ( .A(net362232), .B(net362231), .Z(net377576) );
  XNOR2_X2 U8637 ( .A(net362232), .B(net362231), .ZN(net362141) );
  INV_X4 U8638 ( .A(net377080), .ZN(net377081) );
  AND3_X4 U8639 ( .A1(net377695), .A2(net362179), .A3(net361984), .ZN(
        net362172) );
  INV_X4 U8640 ( .A(net362257), .ZN(n5839) );
  OAI21_X2 U8641 ( .B1(net362224), .B2(n5839), .A(net368201), .ZN(net362211)
         );
  NAND3_X2 U8642 ( .A1(n5839), .A2(net362255), .A3(net362256), .ZN(net362246)
         );
  INV_X4 U8643 ( .A(n5844), .ZN(n5843) );
  NAND2_X2 U8644 ( .A1(n5843), .A2(net362224), .ZN(net377531) );
  NAND2_X4 U8645 ( .A1(n5843), .A2(net362224), .ZN(net361670) );
  NAND3_X2 U8646 ( .A1(net377909), .A2(net362281), .A3(n5311), .ZN(n5844) );
  NAND2_X4 U8647 ( .A1(net362281), .A2(n5311), .ZN(net362362) );
  NAND3_X4 U8648 ( .A1(net377909), .A2(n5311), .A3(net362281), .ZN(net345751)
         );
  NAND3_X4 U8649 ( .A1(net369137), .A2(n5311), .A3(net362281), .ZN(net362337)
         );
  INV_X32 U8650 ( .A(net368498), .ZN(net362224) );
  INV_X32 U8651 ( .A(net368497), .ZN(net368498) );
  INV_X16 U8652 ( .A(net351631), .ZN(net368497) );
  NAND3_X4 U8653 ( .A1(net364871), .A2(net364870), .A3(n5845), .ZN(net351631)
         );
  NAND3_X4 U8654 ( .A1(net364875), .A2(net364874), .A3(n5846), .ZN(n5845) );
  OAI22_X4 U8655 ( .A1(n5848), .A2(n5847), .B1(net369197), .B2(n5849), .ZN(
        net361263) );
  AOI21_X4 U8656 ( .B1(n5850), .B2(n5851), .A(n5852), .ZN(n5849) );
  INV_X4 U8657 ( .A(net359923), .ZN(n5852) );
  XNOR2_X2 U8658 ( .A(net361295), .B(n5857), .ZN(n5851) );
  BUF_X8 U8659 ( .A(net361292), .Z(n5857) );
  NAND3_X1 U8660 ( .A1(net377501), .A2(n5857), .A3(net361293), .ZN(net361289)
         );
  NAND2_X2 U8661 ( .A1(net361291), .A2(n5857), .ZN(net361290) );
  OAI21_X4 U8662 ( .B1(net361809), .B2(net361291), .A(n5857), .ZN(net361740)
         );
  INV_X4 U8663 ( .A(net361296), .ZN(n5850) );
  NAND2_X2 U8664 ( .A1(n5855), .A2(net361709), .ZN(n5847) );
  XNOR2_X2 U8665 ( .A(n5856), .B(aluBoi_multBoi_temppp[39]), .ZN(n5855) );
  XNOR2_X2 U8666 ( .A(n5856), .B(n5585), .ZN(net359792) );
  OAI21_X4 U8667 ( .B1(n5853), .B2(n5854), .A(n5858), .ZN(n5848) );
  NAND2_X2 U8668 ( .A1(n5860), .A2(n5861), .ZN(n5858) );
  NAND2_X2 U8669 ( .A1(n5859), .A2(aluBoi_multBoi_temppp[41]), .ZN(n5861) );
  INV_X4 U8670 ( .A(net361306), .ZN(n5854) );
  AOI21_X4 U8671 ( .B1(net361307), .B2(net361308), .A(net361309), .ZN(n5853)
         );
  INV_X4 U8672 ( .A(net361029), .ZN(net361025) );
  NAND3_X2 U8673 ( .A1(net361002), .A2(n5863), .A3(net361025), .ZN(net361023)
         );
  BUF_X4 U8674 ( .A(net361022), .Z(n5863) );
  OAI21_X2 U8675 ( .B1(net361020), .B2(net361021), .A(n5863), .ZN(net361018)
         );
  INV_X8 U8676 ( .A(net360926), .ZN(net360618) );
  NAND2_X4 U8677 ( .A1(net360617), .A2(net360618), .ZN(net360299) );
  NAND2_X4 U8678 ( .A1(net360617), .A2(net360618), .ZN(net360651) );
  INV_X4 U8679 ( .A(net361030), .ZN(n5862) );
  NAND4_X2 U8680 ( .A1(net361834), .A2(net361833), .A3(net361828), .A4(
        net361835), .ZN(net361356) );
  INV_X4 U8681 ( .A(net362112), .ZN(net378432) );
  INV_X8 U8682 ( .A(net362113), .ZN(net362112) );
  NOR2_X2 U8683 ( .A1(net377355), .A2(net362112), .ZN(net362109) );
  NOR2_X2 U8684 ( .A1(net362112), .A2(net377355), .ZN(net362122) );
  NAND2_X4 U8685 ( .A1(net376960), .A2(net376961), .ZN(net377530) );
  XNOR2_X2 U8686 ( .A(net362117), .B(n10748), .ZN(net362097) );
  INV_X1 U8687 ( .A(net359504), .ZN(net369096) );
  OAI21_X1 U8688 ( .B1(net359504), .B2(net359762), .A(net100619), .ZN(
        net359761) );
  INV_X2 U8689 ( .A(net360017), .ZN(net360014) );
  OAI21_X2 U8690 ( .B1(net359678), .B2(n5864), .A(n5865), .ZN(net360015) );
  NAND2_X1 U8691 ( .A1(net359520), .A2(net359905), .ZN(n5865) );
  AOI21_X4 U8692 ( .B1(net359676), .B2(net377900), .A(net359474), .ZN(
        net360003) );
  INV_X8 U8693 ( .A(net359675), .ZN(net359474) );
  NAND2_X2 U8694 ( .A1(net361411), .A2(net361410), .ZN(net361081) );
  NAND3_X2 U8695 ( .A1(net361073), .A2(n11120), .A3(net369287), .ZN(net361411)
         );
  NAND2_X4 U8696 ( .A1(net362158), .A2(net362159), .ZN(net362051) );
  NAND2_X2 U8697 ( .A1(net362131), .A2(net362051), .ZN(net362149) );
  NAND3_X1 U8698 ( .A1(net362049), .A2(net362050), .A3(net362051), .ZN(
        net362048) );
  INV_X4 U8699 ( .A(net362051), .ZN(net362153) );
  NAND2_X1 U8700 ( .A1(net362317), .A2(net362218), .ZN(net362139) );
  NAND3_X2 U8701 ( .A1(net362063), .A2(net362138), .A3(net362139), .ZN(
        net362131) );
  XNOR2_X2 U8702 ( .A(n5866), .B(net362327), .ZN(net362063) );
  INV_X2 U8703 ( .A(net362063), .ZN(net362062) );
  NAND2_X4 U8704 ( .A1(net375434), .A2(net362330), .ZN(n5866) );
  NAND2_X1 U8705 ( .A1(net362218), .A2(net362318), .ZN(net362138) );
  OAI21_X4 U8706 ( .B1(net368181), .B2(n4981), .A(n5867), .ZN(net361080) );
  NAND2_X2 U8707 ( .A1(net359603), .A2(net368519), .ZN(n5867) );
  INV_X4 U8708 ( .A(net100474), .ZN(net368518) );
  OAI21_X1 U8709 ( .B1(n5868), .B2(n5310), .A(net363049), .ZN(net100474) );
  INV_X4 U8710 ( .A(net363047), .ZN(n5868) );
  INV_X16 U8711 ( .A(net368436), .ZN(net359603) );
  INV_X32 U8712 ( .A(net368435), .ZN(net368436) );
  NOR2_X2 U8713 ( .A1(net359465), .A2(net359474), .ZN(net359473) );
  NOR2_X1 U8714 ( .A1(net359772), .A2(net359512), .ZN(net359770) );
  OAI211_X2 U8715 ( .C1(n12332), .C2(net359515), .A(net359679), .B(net359680), 
        .ZN(net359481) );
  NAND4_X2 U8716 ( .A1(net365032), .A2(net365033), .A3(net365030), .A4(
        net365031), .ZN(net377481) );
  INV_X16 U8717 ( .A(net375650), .ZN(net367041) );
  NAND3_X2 U8718 ( .A1(n11565), .A2(n11563), .A3(n11564), .ZN(n11691) );
  INV_X4 U8719 ( .A(n6785), .ZN(n6492) );
  INV_X8 U8720 ( .A(net376574), .ZN(net378488) );
  INV_X4 U8721 ( .A(n10916), .ZN(n5869) );
  NAND2_X4 U8722 ( .A1(n10670), .A2(n6127), .ZN(n10601) );
  NAND2_X1 U8723 ( .A1(regBoiz_regfile_14__16_), .A2(n6695), .ZN(n967) );
  BUF_X8 U8724 ( .A(n10625), .Z(n5870) );
  NAND3_X1 U8725 ( .A1(n12022), .A2(n12002), .A3(n12023), .ZN(n12103) );
  NAND2_X2 U8726 ( .A1(n11528), .A2(n11609), .ZN(n9899) );
  NAND3_X2 U8727 ( .A1(n11485), .A2(n11530), .A3(n11484), .ZN(n11486) );
  XNOR2_X1 U8728 ( .A(n11529), .B(n6519), .ZN(n11863) );
  NAND2_X2 U8729 ( .A1(n6208), .A2(n11805), .ZN(n11733) );
  NAND4_X4 U8730 ( .A1(n9095), .A2(n9097), .A3(n8718), .A4(n9091), .ZN(n9100)
         );
  NAND2_X2 U8731 ( .A1(n11834), .A2(n12096), .ZN(n6156) );
  INV_X2 U8732 ( .A(net377530), .ZN(n10589) );
  NAND2_X4 U8733 ( .A1(n10834), .A2(n10833), .ZN(n10856) );
  NAND3_X2 U8734 ( .A1(n11057), .A2(n11058), .A3(n11180), .ZN(n5873) );
  NAND3_X2 U8735 ( .A1(n11057), .A2(n11058), .A3(n11180), .ZN(n11254) );
  INV_X2 U8736 ( .A(n12370), .ZN(n5874) );
  INV_X4 U8737 ( .A(n5874), .ZN(n5875) );
  NAND3_X4 U8738 ( .A1(n10746), .A2(n11071), .A3(net368201), .ZN(n10631) );
  NAND2_X4 U8739 ( .A1(net360904), .A2(n6543), .ZN(n10688) );
  NAND2_X2 U8740 ( .A1(n11725), .A2(n9802), .ZN(n9810) );
  INV_X4 U8741 ( .A(n12459), .ZN(n5877) );
  INV_X8 U8742 ( .A(n5877), .ZN(n5878) );
  XNOR2_X2 U8743 ( .A(n8719), .B(n10346), .ZN(n5879) );
  INV_X8 U8744 ( .A(n5879), .ZN(n9091) );
  MUX2_X2 U8745 ( .A(n7577), .B(n7578), .S(net375721), .Z(n7579) );
  INV_X1 U8746 ( .A(n11875), .ZN(n11877) );
  XNOR2_X2 U8747 ( .A(n11847), .B(n11848), .ZN(n5880) );
  NOR2_X4 U8748 ( .A1(net369206), .A2(net366953), .ZN(n5959) );
  INV_X16 U8749 ( .A(net366939), .ZN(net366953) );
  NAND3_X1 U8750 ( .A1(n11472), .A2(n11374), .A3(n11641), .ZN(n11473) );
  NAND3_X2 U8751 ( .A1(net368213), .A2(n10614), .A3(n11071), .ZN(n10615) );
  INV_X4 U8752 ( .A(net359450), .ZN(net359447) );
  NAND2_X4 U8753 ( .A1(n10694), .A2(n10693), .ZN(net378405) );
  NAND2_X4 U8754 ( .A1(net362270), .A2(net362297), .ZN(net362240) );
  INV_X2 U8755 ( .A(n11637), .ZN(n11638) );
  NAND2_X2 U8756 ( .A1(n10855), .A2(n11024), .ZN(n10806) );
  XNOR2_X2 U8757 ( .A(n11864), .B(n5885), .ZN(n5884) );
  XOR2_X2 U8758 ( .A(n11900), .B(n5996), .Z(n5885) );
  NOR2_X4 U8759 ( .A1(n10915), .A2(n10889), .ZN(n10890) );
  NAND2_X1 U8760 ( .A1(regBoiz_regfile_24__28_), .A2(n6734), .ZN(n585) );
  NOR2_X4 U8761 ( .A1(n5520), .A2(n12666), .ZN(n5886) );
  INV_X4 U8762 ( .A(n5886), .ZN(n12660) );
  NAND2_X4 U8763 ( .A1(iaddr[25]), .A2(n12667), .ZN(n12666) );
  XNOR2_X2 U8764 ( .A(n11154), .B(n6427), .ZN(n11151) );
  NAND2_X4 U8765 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  XNOR2_X1 U8766 ( .A(n10887), .B(n6539), .ZN(n5974) );
  AOI211_X2 U8767 ( .C1(n11014), .C2(n11389), .A(n11013), .B(n11012), .ZN(
        n11015) );
  NOR2_X2 U8768 ( .A1(n10985), .A2(n11014), .ZN(n10986) );
  NAND2_X4 U8769 ( .A1(n6010), .A2(n10548), .ZN(n10518) );
  INV_X2 U8770 ( .A(n11556), .ZN(n5887) );
  OAI21_X2 U8771 ( .B1(n12056), .B2(n5001), .A(n6509), .ZN(n12058) );
  INV_X8 U8772 ( .A(net361015), .ZN(net361013) );
  NAND2_X4 U8773 ( .A1(n11416), .A2(n11417), .ZN(n11734) );
  NOR2_X4 U8774 ( .A1(n6431), .A2(n12292), .ZN(n12101) );
  XNOR2_X2 U8775 ( .A(n5889), .B(n10793), .ZN(n10833) );
  NAND2_X4 U8776 ( .A1(n12531), .A2(n12530), .ZN(net359676) );
  INV_X1 U8777 ( .A(n12357), .ZN(n12197) );
  NOR2_X2 U8778 ( .A1(n12429), .A2(n12471), .ZN(n12430) );
  INV_X2 U8779 ( .A(n12471), .ZN(n12362) );
  NOR2_X2 U8780 ( .A1(n5926), .A2(n12471), .ZN(n12363) );
  INV_X8 U8781 ( .A(n10989), .ZN(n10984) );
  INV_X8 U8782 ( .A(n10543), .ZN(n10582) );
  OAI22_X4 U8783 ( .A1(n11764), .A2(net368467), .B1(n12020), .B2(net368211), 
        .ZN(n5890) );
  NAND3_X2 U8784 ( .A1(n11611), .A2(n11610), .A3(n11609), .ZN(n5891) );
  NAND2_X2 U8785 ( .A1(n10563), .A2(n10562), .ZN(n13523) );
  OAI21_X2 U8786 ( .B1(net368185), .B2(n10752), .A(n10747), .ZN(n11021) );
  NAND2_X4 U8787 ( .A1(n10509), .A2(n10526), .ZN(n10520) );
  NAND2_X4 U8788 ( .A1(n11234), .A2(n11312), .ZN(n11241) );
  NAND2_X1 U8789 ( .A1(n12030), .A2(n12093), .ZN(n12099) );
  INV_X16 U8790 ( .A(n11552), .ZN(n5893) );
  OAI21_X2 U8791 ( .B1(n10529), .B2(n10530), .A(net368201), .ZN(n10531) );
  NAND2_X4 U8792 ( .A1(n11299), .A2(n6525), .ZN(n5896) );
  OAI22_X4 U8793 ( .A1(net362216), .A2(net362141), .B1(n6130), .B2(n10542), 
        .ZN(n10543) );
  NAND2_X1 U8794 ( .A1(net361512), .A2(n10989), .ZN(n10945) );
  XNOR2_X2 U8795 ( .A(net361713), .B(net361291), .ZN(net378052) );
  INV_X2 U8796 ( .A(net361713), .ZN(net361809) );
  NOR2_X2 U8797 ( .A1(net376602), .A2(net377531), .ZN(n10550) );
  INV_X4 U8798 ( .A(n5897), .ZN(n5898) );
  NAND2_X4 U8799 ( .A1(n11118), .A2(n11117), .ZN(n11082) );
  AOI21_X4 U8800 ( .B1(n11020), .B2(net361372), .A(n11019), .ZN(n11081) );
  INV_X16 U8801 ( .A(net369232), .ZN(net378318) );
  INV_X2 U8802 ( .A(n10610), .ZN(n5899) );
  NOR3_X4 U8803 ( .A1(n5987), .A2(n6527), .A3(n6194), .ZN(n11297) );
  NAND4_X4 U8804 ( .A1(n8073), .A2(n6008), .A3(n6787), .A4(net375876), .ZN(
        n10453) );
  NAND4_X2 U8805 ( .A1(n8073), .A2(n6008), .A3(n6787), .A4(net375876), .ZN(
        n6075) );
  MUX2_X2 U8806 ( .A(n7513), .B(n7512), .S(net366933), .Z(n5900) );
  MUX2_X2 U8807 ( .A(n7511), .B(n7510), .S(net366969), .Z(n7512) );
  NAND2_X2 U8808 ( .A1(net368215), .A2(n11000), .ZN(n10706) );
  NAND2_X2 U8809 ( .A1(n10505), .A2(n10563), .ZN(n10506) );
  XOR2_X1 U8810 ( .A(n10734), .B(n10733), .Z(n5901) );
  NAND2_X4 U8811 ( .A1(n10789), .A2(n10790), .ZN(n10734) );
  INV_X1 U8812 ( .A(n10554), .ZN(n5902) );
  INV_X8 U8813 ( .A(n10551), .ZN(n10554) );
  XNOR2_X2 U8814 ( .A(n5904), .B(n12281), .ZN(n5903) );
  XOR2_X2 U8815 ( .A(n12382), .B(n12469), .Z(n5904) );
  AOI22_X4 U8816 ( .A1(n11025), .A2(n11024), .B1(n11023), .B2(n11024), .ZN(
        net361541) );
  OAI21_X1 U8817 ( .B1(net362125), .B2(net362126), .A(net362091), .ZN(n10598)
         );
  XNOR2_X1 U8818 ( .A(n6427), .B(n10854), .ZN(n5905) );
  MUX2_X2 U8819 ( .A(n7525), .B(n7524), .S(net366971), .Z(n7526) );
  INV_X4 U8820 ( .A(n12415), .ZN(n12405) );
  NAND2_X4 U8821 ( .A1(n11813), .A2(n11814), .ZN(n11820) );
  OAI22_X4 U8822 ( .A1(net360490), .A2(net368467), .B1(net360206), .B2(
        net368211), .ZN(n11813) );
  OAI211_X4 U8823 ( .C1(n7806), .C2(n7805), .A(net361491), .B(n7804), .ZN(
        n5907) );
  NAND3_X2 U8824 ( .A1(n12354), .A2(n12460), .A3(n12353), .ZN(n12355) );
  OAI21_X2 U8825 ( .B1(n10589), .B2(net361913), .A(net378060), .ZN(net362142)
         );
  NAND2_X4 U8826 ( .A1(net360821), .A2(n6543), .ZN(n10616) );
  INV_X16 U8827 ( .A(n6542), .ZN(n6543) );
  INV_X2 U8828 ( .A(n12376), .ZN(n5908) );
  INV_X4 U8829 ( .A(n5908), .ZN(n5909) );
  INV_X2 U8830 ( .A(n10760), .ZN(n5910) );
  INV_X4 U8831 ( .A(n10859), .ZN(n10760) );
  INV_X2 U8832 ( .A(n10837), .ZN(n10823) );
  NOR2_X4 U8833 ( .A1(n12169), .A2(n12171), .ZN(n5911) );
  INV_X4 U8834 ( .A(n5911), .ZN(n12070) );
  NAND2_X2 U8835 ( .A1(n11984), .A2(n11983), .ZN(n12168) );
  INV_X8 U8836 ( .A(n6425), .ZN(n11402) );
  XNOR2_X2 U8837 ( .A(net362094), .B(net362095), .ZN(n5912) );
  XNOR2_X1 U8838 ( .A(net362094), .B(net362095), .ZN(n5913) );
  INV_X1 U8839 ( .A(n12172), .ZN(n5914) );
  AOI22_X4 U8840 ( .A1(n5916), .A2(idOut_110_), .B1(n5917), .B2(n5918), .ZN(
        n5915) );
  NOR2_X2 U8841 ( .A1(n11742), .A2(n11736), .ZN(n11737) );
  OAI21_X4 U8842 ( .B1(n11141), .B2(net361361), .A(n5985), .ZN(n11361) );
  INV_X4 U8843 ( .A(n11339), .ZN(n5985) );
  NAND2_X4 U8844 ( .A1(n12400), .A2(n12401), .ZN(n12403) );
  XNOR2_X2 U8845 ( .A(n11788), .B(n5920), .ZN(n5919) );
  INV_X4 U8846 ( .A(n5919), .ZN(n11868) );
  INV_X4 U8847 ( .A(net362052), .ZN(net362047) );
  AOI21_X4 U8848 ( .B1(n11082), .B2(net369286), .A(n11026), .ZN(n11020) );
  NAND3_X4 U8849 ( .A1(n11547), .A2(n11342), .A3(n11324), .ZN(n11367) );
  NAND2_X4 U8850 ( .A1(n10532), .A2(n10533), .ZN(net362231) );
  INV_X8 U8851 ( .A(net375642), .ZN(net376076) );
  NAND2_X4 U8852 ( .A1(n11923), .A2(n11932), .ZN(n11924) );
  NOR2_X4 U8853 ( .A1(n13533), .A2(n6535), .ZN(n5922) );
  INV_X2 U8854 ( .A(n11736), .ZN(n5923) );
  AOI21_X4 U8855 ( .B1(n6089), .B2(n10874), .A(n10864), .ZN(n10865) );
  XNOR2_X2 U8856 ( .A(n11336), .B(n11337), .ZN(n5924) );
  INV_X4 U8857 ( .A(n11336), .ZN(n11161) );
  NAND4_X2 U8858 ( .A1(n11927), .A2(n11925), .A3(n11926), .A4(n11924), .ZN(
        n5925) );
  NAND4_X2 U8859 ( .A1(n11927), .A2(n11925), .A3(n11926), .A4(n11924), .ZN(
        n11941) );
  NAND4_X2 U8860 ( .A1(n12255), .A2(n12256), .A3(n12257), .A4(n12568), .ZN(
        n12262) );
  CLKBUF_X3 U8861 ( .A(n12463), .Z(n5926) );
  NAND2_X4 U8862 ( .A1(net375713), .A2(n7803), .ZN(n7804) );
  NAND2_X4 U8863 ( .A1(n11559), .A2(n11558), .ZN(n11657) );
  OAI21_X1 U8864 ( .B1(n6553), .B2(n11475), .A(n5893), .ZN(n5928) );
  INV_X8 U8865 ( .A(n11797), .ZN(n11475) );
  XNOR2_X2 U8866 ( .A(n11346), .B(n5923), .ZN(n11332) );
  INV_X4 U8867 ( .A(n11346), .ZN(n11330) );
  INV_X8 U8868 ( .A(n11597), .ZN(n11627) );
  NOR3_X2 U8869 ( .A1(n12003), .A2(n12078), .A3(n12274), .ZN(n12008) );
  NOR3_X2 U8870 ( .A1(n12464), .A2(n12003), .A3(n12274), .ZN(n12007) );
  INV_X4 U8871 ( .A(n12165), .ZN(n12274) );
  NOR2_X4 U8872 ( .A1(n13533), .A2(n6535), .ZN(n5929) );
  INV_X4 U8873 ( .A(n5922), .ZN(n11184) );
  NAND2_X4 U8874 ( .A1(n11774), .A2(n12055), .ZN(net360206) );
  NOR3_X4 U8875 ( .A1(n10912), .A2(n10913), .A3(n6539), .ZN(n10928) );
  MUX2_X2 U8876 ( .A(n5931), .B(n5932), .S(net376077), .Z(n5930) );
  INV_X4 U8877 ( .A(n11898), .ZN(n5933) );
  AND2_X4 U8878 ( .A1(n6109), .A2(n6110), .ZN(n7562) );
  OAI21_X4 U8879 ( .B1(n10767), .B2(n10766), .A(n10765), .ZN(n11166) );
  INV_X4 U8880 ( .A(n12136), .ZN(n5934) );
  NAND2_X4 U8881 ( .A1(n12028), .A2(n12079), .ZN(n11834) );
  INV_X2 U8882 ( .A(n11361), .ZN(n11158) );
  NOR2_X4 U8883 ( .A1(n6059), .A2(n12119), .ZN(n11566) );
  INV_X8 U8884 ( .A(n12450), .ZN(n5937) );
  INV_X8 U8885 ( .A(n12448), .ZN(n12450) );
  AND3_X4 U8886 ( .A1(n11945), .A2(n11920), .A3(n11963), .ZN(n11936) );
  OAI21_X1 U8887 ( .B1(n12560), .B2(n12390), .A(n12559), .ZN(n12589) );
  INV_X8 U8888 ( .A(n12271), .ZN(n12358) );
  INV_X1 U8889 ( .A(net360617), .ZN(net377462) );
  INV_X8 U8890 ( .A(n11375), .ZN(n5938) );
  INV_X16 U8891 ( .A(n5938), .ZN(n5939) );
  INV_X4 U8892 ( .A(n12404), .ZN(n12414) );
  NAND2_X4 U8893 ( .A1(n12392), .A2(n12375), .ZN(n12404) );
  NAND2_X2 U8894 ( .A1(n12405), .A2(n12407), .ZN(n12387) );
  INV_X4 U8895 ( .A(net361748), .ZN(net376121) );
  INV_X4 U8896 ( .A(regBoiz_N15), .ZN(net378137) );
  INV_X8 U8897 ( .A(net378137), .ZN(net378138) );
  INV_X4 U8898 ( .A(n5940), .ZN(ifInst[1]) );
  INV_X8 U8899 ( .A(n11153), .ZN(n11337) );
  NOR3_X2 U8900 ( .A1(n12162), .A2(n6124), .A3(n5989), .ZN(n12196) );
  INV_X4 U8901 ( .A(net361509), .ZN(net378128) );
  INV_X8 U8902 ( .A(n11988), .ZN(n5943) );
  INV_X8 U8903 ( .A(n12190), .ZN(n11988) );
  OAI22_X4 U8904 ( .A1(net360713), .A2(net368467), .B1(net377575), .B2(
        net368211), .ZN(n11716) );
  XNOR2_X2 U8905 ( .A(aluRw[4]), .B(n6783), .ZN(n6995) );
  INV_X1 U8906 ( .A(net369197), .ZN(net375948) );
  INV_X2 U8907 ( .A(n11305), .ZN(n5946) );
  NAND3_X2 U8908 ( .A1(n8120), .A2(n8119), .A3(net368781), .ZN(net364874) );
  INV_X4 U8909 ( .A(n10849), .ZN(n5947) );
  NOR2_X4 U8910 ( .A1(n9817), .A2(n9816), .ZN(n5948) );
  NAND2_X4 U8911 ( .A1(n11664), .A2(n11691), .ZN(n11913) );
  OAI21_X4 U8912 ( .B1(n11546), .B2(net368195), .A(n11461), .ZN(n11463) );
  XNOR2_X2 U8913 ( .A(n5949), .B(net376642), .ZN(n6997) );
  NOR2_X2 U8914 ( .A1(n5989), .A2(n12436), .ZN(n12198) );
  NAND2_X2 U8915 ( .A1(n11001), .A2(n11197), .ZN(n11002) );
  INV_X2 U8916 ( .A(n6194), .ZN(n11197) );
  XNOR2_X2 U8917 ( .A(n5905), .B(n11154), .ZN(n5950) );
  XNOR2_X1 U8918 ( .A(n10627), .B(n10577), .ZN(n5951) );
  NAND3_X2 U8919 ( .A1(n5881), .A2(n10634), .A3(n10635), .ZN(n10577) );
  OAI21_X4 U8920 ( .B1(n10510), .B2(net377937), .A(net362297), .ZN(n5952) );
  NAND2_X1 U8921 ( .A1(n9065), .A2(n9064), .ZN(n9466) );
  NOR2_X2 U8922 ( .A1(n9074), .A2(n9073), .ZN(n9077) );
  NOR3_X1 U8923 ( .A1(n9066), .A2(n9104), .A3(n9073), .ZN(n9069) );
  INV_X4 U8924 ( .A(n4993), .ZN(n10991) );
  OAI21_X4 U8925 ( .B1(n5332), .B2(n11006), .A(n11005), .ZN(n5953) );
  NAND3_X4 U8926 ( .A1(n5881), .A2(n10635), .A3(n10634), .ZN(n10639) );
  INV_X4 U8927 ( .A(n6100), .ZN(n11740) );
  NOR2_X4 U8928 ( .A1(n5955), .A2(n10500), .ZN(n5954) );
  INV_X4 U8929 ( .A(n5954), .ZN(n9080) );
  INV_X2 U8930 ( .A(n13140), .ZN(n13141) );
  NAND2_X1 U8931 ( .A1(n13140), .A2(n13129), .ZN(n9046) );
  INV_X2 U8932 ( .A(n9784), .ZN(n5956) );
  INV_X2 U8933 ( .A(n10513), .ZN(n9784) );
  INV_X8 U8934 ( .A(n8879), .ZN(n9095) );
  INV_X1 U8935 ( .A(n12361), .ZN(n5957) );
  INV_X4 U8936 ( .A(n11229), .ZN(n5987) );
  OAI22_X4 U8937 ( .A1(n10998), .A2(net368462), .B1(n11331), .B2(net368195), 
        .ZN(n5958) );
  OAI22_X2 U8938 ( .A1(n10998), .A2(net368462), .B1(n11331), .B2(net368195), 
        .ZN(n11457) );
  NOR2_X1 U8939 ( .A1(n9095), .A2(n9087), .ZN(n9090) );
  NAND2_X2 U8940 ( .A1(net361293), .A2(n11166), .ZN(net361713) );
  NAND2_X4 U8941 ( .A1(n11600), .A2(n11599), .ZN(n11602) );
  NAND2_X4 U8942 ( .A1(net375434), .A2(net362330), .ZN(n10486) );
  NAND2_X4 U8943 ( .A1(n5907), .A2(n10703), .ZN(n10724) );
  NAND2_X4 U8944 ( .A1(n10704), .A2(n10703), .ZN(n10770) );
  INV_X1 U8945 ( .A(n11847), .ZN(n11761) );
  NAND2_X2 U8946 ( .A1(net369200), .A2(net375717), .ZN(n5960) );
  NAND2_X4 U8947 ( .A1(net369200), .A2(net375717), .ZN(n5961) );
  XNOR2_X2 U8948 ( .A(n11079), .B(n11204), .ZN(n5962) );
  OAI21_X1 U8949 ( .B1(n8112), .B2(n8111), .A(net366967), .ZN(n8120) );
  OAI21_X1 U8950 ( .B1(n8118), .B2(n8117), .A(net366999), .ZN(n8119) );
  NOR2_X1 U8951 ( .A1(n6553), .A2(n6432), .ZN(n11710) );
  XNOR2_X2 U8952 ( .A(n11638), .B(n11583), .ZN(n5963) );
  INV_X4 U8953 ( .A(n5963), .ZN(n11750) );
  INV_X2 U8954 ( .A(n11022), .ZN(n11023) );
  NOR2_X4 U8955 ( .A1(n11626), .A2(n11388), .ZN(n5964) );
  INV_X2 U8956 ( .A(n11626), .ZN(n11598) );
  NAND2_X4 U8957 ( .A1(n11593), .A2(n11646), .ZN(n11626) );
  INV_X8 U8958 ( .A(n11458), .ZN(n11388) );
  INV_X1 U8959 ( .A(n10660), .ZN(n10659) );
  NAND2_X4 U8960 ( .A1(n11291), .A2(n11292), .ZN(n11250) );
  XNOR2_X2 U8961 ( .A(n10795), .B(net361548), .ZN(n5965) );
  INV_X8 U8962 ( .A(net369210), .ZN(net375727) );
  BUF_X4 U8963 ( .A(net361886), .Z(net378013) );
  OAI21_X4 U8964 ( .B1(n12424), .B2(n5027), .A(n12422), .ZN(n12457) );
  NAND2_X1 U8965 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  NAND2_X4 U8966 ( .A1(n11402), .A2(n11401), .ZN(n11390) );
  OAI21_X2 U8967 ( .B1(n5682), .B2(n6769), .A(n181), .ZN(n4429) );
  INV_X16 U8968 ( .A(n13521), .ZN(n6526) );
  INV_X1 U8969 ( .A(n12437), .ZN(n5968) );
  INV_X2 U8970 ( .A(n5968), .ZN(n5969) );
  XNOR2_X2 U8971 ( .A(net361547), .B(net361629), .ZN(n10795) );
  INV_X8 U8972 ( .A(net361546), .ZN(net361547) );
  XNOR2_X2 U8973 ( .A(n10980), .B(n10979), .ZN(n5970) );
  INV_X1 U8974 ( .A(n6535), .ZN(n11041) );
  XNOR2_X1 U8975 ( .A(n11003), .B(n8450), .ZN(n9470) );
  AOI21_X2 U8976 ( .B1(n9657), .B2(n6560), .A(n11003), .ZN(n9658) );
  NAND3_X2 U8977 ( .A1(n8937), .A2(n8930), .A3(n8936), .ZN(n8931) );
  NOR2_X1 U8978 ( .A1(n10895), .A2(n10894), .ZN(n10896) );
  INV_X2 U8979 ( .A(n11869), .ZN(n11874) );
  NAND3_X2 U8980 ( .A1(net366919), .A2(net369316), .A3(n6782), .ZN(n7976) );
  NAND3_X2 U8981 ( .A1(n6782), .A2(net366947), .A3(net369316), .ZN(n9854) );
  NOR2_X2 U8982 ( .A1(net369316), .A2(n6782), .ZN(n11051) );
  AOI21_X2 U8983 ( .B1(regBoiz_regfile_24__30_), .B2(n6782), .A(net366925), 
        .ZN(n8079) );
  AOI21_X2 U8984 ( .B1(regBoiz_regfile_26__30_), .B2(n6782), .A(net366925), 
        .ZN(n8076) );
  NOR2_X2 U8985 ( .A1(n6782), .A2(n5576), .ZN(n8133) );
  NOR2_X2 U8986 ( .A1(n6782), .A2(n5577), .ZN(n8137) );
  NAND4_X2 U8987 ( .A1(n11055), .A2(net361491), .A3(n11056), .A4(n6787), .ZN(
        n11057) );
  OAI21_X2 U8988 ( .B1(n5692), .B2(n7699), .A(n6793), .ZN(n7703) );
  INV_X8 U8989 ( .A(n6796), .ZN(n6793) );
  OAI21_X2 U8990 ( .B1(n7684), .B2(n7683), .A(n6794), .ZN(n7688) );
  NAND3_X1 U8991 ( .A1(n7332), .A2(n6794), .A3(net366953), .ZN(n7333) );
  NAND2_X1 U8992 ( .A1(regBoiz_regfile_11__30_), .A2(n6794), .ZN(n8110) );
  NAND2_X1 U8993 ( .A1(regBoiz_regfile_2__30_), .A2(n6794), .ZN(n8098) );
  NAND2_X1 U8994 ( .A1(regBoiz_regfile_0__30_), .A2(n6794), .ZN(n8092) );
  AOI21_X2 U8995 ( .B1(regBoiz_regfile_7__31_), .B2(n6793), .A(net366951), 
        .ZN(n8145) );
  AOI21_X1 U8996 ( .B1(regBoiz_regfile_5__31_), .B2(n6793), .A(net366951), 
        .ZN(n8142) );
  AOI21_X2 U8997 ( .B1(regBoiz_regfile_24__19_), .B2(net366949), .A(n6793), 
        .ZN(n7628) );
  OAI21_X2 U8998 ( .B1(n5694), .B2(n7678), .A(n6793), .ZN(n7681) );
  OAI21_X2 U8999 ( .B1(n5695), .B2(n7689), .A(n6793), .ZN(n7695) );
  OAI21_X2 U9000 ( .B1(n5693), .B2(n7720), .A(n6793), .ZN(n7725) );
  OAI21_X4 U9001 ( .B1(n9892), .B2(n10697), .A(n11192), .ZN(n9893) );
  INV_X2 U9002 ( .A(n12256), .ZN(n5971) );
  XNOR2_X2 U9003 ( .A(n9677), .B(n10415), .ZN(n8587) );
  INV_X2 U9004 ( .A(n10415), .ZN(n9631) );
  NAND3_X2 U9005 ( .A1(n8585), .A2(n8584), .A3(n8583), .ZN(n10415) );
  NAND4_X2 U9006 ( .A1(n12123), .A2(n11934), .A3(n12122), .A4(net360297), .ZN(
        n11935) );
  OAI21_X2 U9007 ( .B1(n8183), .B2(n8182), .A(n8181), .ZN(n10513) );
  INV_X1 U9008 ( .A(net368584), .ZN(net360490) );
  XNOR2_X2 U9009 ( .A(n5045), .B(n11943), .ZN(net360261) );
  INV_X1 U9010 ( .A(n11741), .ZN(n5973) );
  OAI21_X4 U9011 ( .B1(n10767), .B2(n10766), .A(n10765), .ZN(net377501) );
  OAI21_X1 U9012 ( .B1(net361326), .B2(net361274), .A(net361327), .ZN(
        net361321) );
  BUF_X8 U9013 ( .A(n11901), .Z(n5975) );
  OAI211_X2 U9014 ( .C1(n6119), .C2(n11642), .A(n11458), .B(n11641), .ZN(
        n11404) );
  INV_X1 U9015 ( .A(n11660), .ZN(n5976) );
  INV_X8 U9016 ( .A(n11303), .ZN(n11242) );
  NAND2_X4 U9017 ( .A1(n11104), .A2(n11103), .ZN(n11106) );
  OAI21_X4 U9018 ( .B1(n8183), .B2(n8182), .A(n8181), .ZN(net377909) );
  INV_X8 U9019 ( .A(n10955), .ZN(n6435) );
  NOR3_X1 U9020 ( .A1(net359765), .A2(n12518), .A3(net359520), .ZN(n12520) );
  INV_X1 U9021 ( .A(n11310), .ZN(n5979) );
  INV_X2 U9022 ( .A(n5979), .ZN(n5980) );
  NAND2_X2 U9023 ( .A1(net362110), .A2(net361913), .ZN(n10590) );
  NAND2_X2 U9024 ( .A1(n10591), .A2(n10590), .ZN(net362117) );
  NAND2_X1 U9025 ( .A1(n12153), .A2(n12406), .ZN(n12378) );
  NOR2_X4 U9026 ( .A1(n12420), .A2(n12421), .ZN(n12424) );
  XNOR2_X2 U9027 ( .A(n11990), .B(n6096), .ZN(n5982) );
  INV_X4 U9028 ( .A(n6096), .ZN(n6097) );
  INV_X2 U9029 ( .A(n4977), .ZN(n6096) );
  INV_X8 U9030 ( .A(n10703), .ZN(n9883) );
  INV_X4 U9031 ( .A(n5332), .ZN(n5983) );
  NAND2_X4 U9032 ( .A1(n9878), .A2(n6788), .ZN(n6174) );
  OAI21_X2 U9033 ( .B1(n5651), .B2(n6693), .A(n971), .ZN(n3876) );
  INV_X8 U9034 ( .A(n12120), .ZN(n11836) );
  INV_X2 U9035 ( .A(net360235), .ZN(net360297) );
  NAND3_X1 U9036 ( .A1(net366907), .A2(net366919), .A3(net366997), .ZN(n8003)
         );
  INV_X4 U9037 ( .A(n6351), .ZN(n7107) );
  INV_X1 U9038 ( .A(n11544), .ZN(n6151) );
  NAND2_X4 U9039 ( .A1(n5890), .A2(n11780), .ZN(n11786) );
  INV_X2 U9040 ( .A(n12243), .ZN(n12153) );
  OAI21_X4 U9041 ( .B1(n11190), .B2(n11191), .A(n11189), .ZN(n11218) );
  NOR3_X4 U9042 ( .A1(n11186), .A2(n5987), .A3(n6194), .ZN(n11190) );
  INV_X16 U9043 ( .A(n6250), .ZN(n6251) );
  INV_X4 U9044 ( .A(n11676), .ZN(n5986) );
  INV_X2 U9045 ( .A(n11675), .ZN(n11676) );
  AOI21_X2 U9046 ( .B1(n6427), .B2(n6071), .A(n11152), .ZN(n11038) );
  XNOR2_X2 U9047 ( .A(n12403), .B(n6212), .ZN(n5988) );
  AOI21_X2 U9048 ( .B1(n5553), .B2(n7592), .A(net365399), .ZN(n7593) );
  MUX2_X2 U9049 ( .A(n7591), .B(n7590), .S(net366971), .Z(n7592) );
  OAI21_X1 U9050 ( .B1(n11311), .B2(n5980), .A(n6529), .ZN(n11313) );
  INV_X8 U9051 ( .A(n12358), .ZN(n5989) );
  INV_X1 U9052 ( .A(n10878), .ZN(n10879) );
  NOR2_X1 U9053 ( .A1(n11329), .A2(n11496), .ZN(n5990) );
  INV_X8 U9054 ( .A(n11409), .ZN(n11496) );
  INV_X8 U9055 ( .A(n10985), .ZN(n6029) );
  NAND2_X4 U9056 ( .A1(n11397), .A2(n5040), .ZN(n11095) );
  INV_X8 U9057 ( .A(n10888), .ZN(n5991) );
  INV_X8 U9058 ( .A(n11096), .ZN(n10888) );
  INV_X2 U9059 ( .A(n11508), .ZN(n11511) );
  NAND2_X4 U9060 ( .A1(n10937), .A2(n6029), .ZN(n11094) );
  NOR2_X2 U9061 ( .A1(n6059), .A2(net360235), .ZN(n11961) );
  NOR3_X2 U9062 ( .A1(n11952), .A2(n11951), .A3(net360235), .ZN(n11956) );
  NAND2_X2 U9063 ( .A1(n11258), .A2(n11736), .ZN(n11260) );
  XNOR2_X2 U9064 ( .A(aluRw[0]), .B(net376222), .ZN(n6996) );
  NAND2_X1 U9065 ( .A1(regBoiz_regfile_27__17_), .A2(n6745), .ZN(n497) );
  NAND4_X2 U9066 ( .A1(n6374), .A2(n11770), .A3(n11729), .A4(n11728), .ZN(
        n5992) );
  NAND4_X2 U9067 ( .A1(n6374), .A2(n11770), .A3(n11729), .A4(n11728), .ZN(
        n11765) );
  XNOR2_X1 U9068 ( .A(n12398), .B(n6113), .ZN(n6065) );
  XNOR2_X2 U9069 ( .A(n11733), .B(n11732), .ZN(n5995) );
  XNOR2_X2 U9070 ( .A(n11733), .B(n11732), .ZN(n5996) );
  NAND2_X2 U9071 ( .A1(n6151), .A2(n11533), .ZN(n6153) );
  AOI21_X1 U9072 ( .B1(n11283), .B2(n11400), .A(n11264), .ZN(n11227) );
  NAND2_X1 U9073 ( .A1(n11283), .A2(n5939), .ZN(n11286) );
  NOR3_X2 U9074 ( .A1(n11228), .A2(n11227), .A3(n5938), .ZN(n11257) );
  INV_X2 U9075 ( .A(n11207), .ZN(n11209) );
  NAND2_X2 U9076 ( .A1(n6427), .A2(n6071), .ZN(n11107) );
  INV_X4 U9077 ( .A(n6367), .ZN(n7800) );
  NAND2_X4 U9078 ( .A1(n11164), .A2(n6009), .ZN(net361319) );
  INV_X8 U9079 ( .A(n12108), .ZN(n12029) );
  INV_X2 U9080 ( .A(net362178), .ZN(net362177) );
  XNOR2_X1 U9081 ( .A(n11855), .B(n11892), .ZN(n11562) );
  INV_X1 U9082 ( .A(n11253), .ZN(n5998) );
  INV_X4 U9083 ( .A(n11470), .ZN(n11253) );
  INV_X4 U9084 ( .A(n6068), .ZN(n12246) );
  INV_X4 U9085 ( .A(n10800), .ZN(n6134) );
  OAI21_X2 U9086 ( .B1(net359673), .B2(n12399), .A(net359675), .ZN(n12484) );
  INV_X2 U9087 ( .A(n12484), .ZN(n12417) );
  AND2_X2 U9088 ( .A1(n11329), .A2(n11408), .ZN(n5999) );
  INV_X8 U9089 ( .A(n11089), .ZN(n11329) );
  INV_X2 U9090 ( .A(net359532), .ZN(net359531) );
  XNOR2_X1 U9091 ( .A(net377947), .B(n5573), .ZN(n12327) );
  AND3_X4 U9092 ( .A1(n11441), .A2(n11500), .A3(n11440), .ZN(n6000) );
  INV_X8 U9093 ( .A(n6000), .ZN(n11738) );
  NAND2_X1 U9094 ( .A1(n12048), .A2(n4994), .ZN(n12174) );
  OAI22_X4 U9095 ( .A1(n11993), .A2(net368467), .B1(n12248), .B2(net368211), 
        .ZN(n12047) );
  AOI21_X4 U9096 ( .B1(n10602), .B2(n10601), .A(n10600), .ZN(n6001) );
  NOR2_X2 U9097 ( .A1(net361547), .A2(net361548), .ZN(net361543) );
  INV_X1 U9098 ( .A(n11792), .ZN(n6002) );
  NAND2_X2 U9099 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  NOR2_X2 U9100 ( .A1(n12524), .A2(net369096), .ZN(n12527) );
  NOR2_X2 U9101 ( .A1(net359761), .A2(n12338), .ZN(n12339) );
  NAND2_X4 U9102 ( .A1(n11893), .A2(n11892), .ZN(n11901) );
  INV_X4 U9103 ( .A(n10918), .ZN(n6003) );
  INV_X4 U9104 ( .A(n12288), .ZN(n6004) );
  INV_X4 U9105 ( .A(n12408), .ZN(n12288) );
  NAND4_X4 U9106 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(net360497), .ZN(
        n11772) );
  INV_X8 U9107 ( .A(n11768), .ZN(n11770) );
  XNOR2_X2 U9108 ( .A(net361906), .B(net377700), .ZN(n6007) );
  AOI21_X4 U9109 ( .B1(n5958), .B2(n5953), .A(n11455), .ZN(n11593) );
  INV_X4 U9110 ( .A(net362177), .ZN(net377695) );
  CLKBUF_X3 U9111 ( .A(net359535), .Z(net377689) );
  INV_X8 U9112 ( .A(n11175), .ZN(n11076) );
  NAND3_X2 U9113 ( .A1(n10438), .A2(n10439), .A3(net375717), .ZN(n6008) );
  INV_X8 U9114 ( .A(n11319), .ZN(n6009) );
  NAND3_X1 U9115 ( .A1(n10512), .A2(n10511), .A3(net361984), .ZN(n6010) );
  NOR2_X4 U9116 ( .A1(n10510), .A2(net377937), .ZN(n10511) );
  XNOR2_X2 U9117 ( .A(n10762), .B(n10763), .ZN(n6011) );
  INV_X4 U9118 ( .A(n6011), .ZN(n10866) );
  NAND3_X1 U9119 ( .A1(net368571), .A2(n11524), .A3(n11523), .ZN(n6012) );
  INV_X4 U9120 ( .A(n11530), .ZN(n11523) );
  INV_X4 U9121 ( .A(n10941), .ZN(n6014) );
  INV_X2 U9122 ( .A(n11115), .ZN(n11141) );
  AOI22_X4 U9123 ( .A1(ifOut_66_), .A2(idBoi_temPC_2_), .B1(n10385), .B2(n9908), .ZN(n10377) );
  OR3_X1 U9124 ( .A1(ifInst[23]), .A2(ifInst[2]), .A3(ifInst[24]), .ZN(n2010)
         );
  NAND4_X1 U9125 ( .A1(n13333), .A2(ifInst[2]), .A3(n5346), .A4(n13288), .ZN(
        n13308) );
  NOR3_X4 U9126 ( .A1(n12385), .A2(n12450), .A3(n12301), .ZN(n6016) );
  INV_X4 U9127 ( .A(n6016), .ZN(n12407) );
  MUX2_X1 U9128 ( .A(n7360), .B(n7359), .S(net366927), .Z(n7361) );
  NAND2_X4 U9129 ( .A1(n10538), .A2(n10545), .ZN(net362158) );
  NAND3_X2 U9130 ( .A1(n10544), .A2(n6194), .A3(net362223), .ZN(n10538) );
  INV_X2 U9131 ( .A(n6017), .ZN(n6018) );
  NAND3_X2 U9132 ( .A1(n12378), .A2(n6004), .A3(n12377), .ZN(n12535) );
  NAND2_X4 U9133 ( .A1(n12245), .A2(n12127), .ZN(n12293) );
  AOI22_X4 U9134 ( .A1(n6036), .A2(n5308), .B1(n5308), .B2(n13280), .ZN(n6019)
         );
  INV_X8 U9135 ( .A(n6019), .ZN(n8712) );
  INV_X8 U9136 ( .A(n9718), .ZN(n6036) );
  NAND3_X2 U9137 ( .A1(n11753), .A2(n11760), .A3(n11752), .ZN(n11871) );
  OAI21_X2 U9138 ( .B1(n5651), .B2(n6697), .A(n937), .ZN(n3877) );
  INV_X2 U9139 ( .A(n6021), .ZN(n6022) );
  AND3_X2 U9140 ( .A1(n10570), .A2(net362322), .A3(n10520), .ZN(n10523) );
  INV_X2 U9141 ( .A(net368498), .ZN(net362322) );
  INV_X4 U9142 ( .A(n11285), .ZN(n6026) );
  INV_X4 U9143 ( .A(n10907), .ZN(n10996) );
  XNOR2_X2 U9144 ( .A(n11483), .B(n11380), .ZN(n11382) );
  NOR2_X1 U9145 ( .A1(n12508), .A2(net359540), .ZN(n12515) );
  NOR2_X4 U9146 ( .A1(n10955), .A2(n10956), .ZN(n10839) );
  NAND2_X4 U9147 ( .A1(n12535), .A2(n12534), .ZN(n12537) );
  XNOR2_X2 U9148 ( .A(n10927), .B(n10987), .ZN(n10983) );
  INV_X8 U9149 ( .A(n11042), .ZN(n10985) );
  NAND2_X4 U9150 ( .A1(n10821), .A2(n5166), .ZN(n11042) );
  NAND3_X2 U9151 ( .A1(n11773), .A2(n11978), .A3(n11977), .ZN(n6027) );
  NOR2_X4 U9152 ( .A1(n4999), .A2(n10912), .ZN(n11066) );
  INV_X16 U9153 ( .A(n11725), .ZN(net377607) );
  NAND3_X2 U9154 ( .A1(n9801), .A2(n9800), .A3(n9799), .ZN(net327826) );
  BUF_X8 U9155 ( .A(n12415), .Z(n6028) );
  XNOR2_X2 U9156 ( .A(n6615), .B(n9677), .ZN(n6055) );
  INV_X2 U9157 ( .A(n6030), .ZN(n6031) );
  NAND3_X2 U9158 ( .A1(n12023), .A2(n12002), .A3(n12022), .ZN(n6032) );
  XNOR2_X2 U9159 ( .A(n12027), .B(n12026), .ZN(n6033) );
  XNOR2_X2 U9160 ( .A(n12464), .B(n12114), .ZN(n12026) );
  OAI211_X2 U9161 ( .C1(n10756), .C2(net361885), .A(net376691), .B(net378013), 
        .ZN(n10757) );
  NOR2_X4 U9162 ( .A1(net361013), .A2(n11361), .ZN(n11362) );
  AOI21_X4 U9163 ( .B1(n11310), .B2(n6529), .A(net368195), .ZN(n11238) );
  XNOR2_X2 U9164 ( .A(n11612), .B(net377607), .ZN(net377575) );
  AOI22_X4 U9165 ( .A1(n6036), .A2(n6037), .B1(n6038), .B2(n13246), .ZN(n6035)
         );
  NAND2_X4 U9166 ( .A1(n11500), .A2(n11646), .ZN(n11501) );
  INV_X4 U9167 ( .A(n10751), .ZN(n6039) );
  INV_X4 U9168 ( .A(n11969), .ZN(n6041) );
  INV_X2 U9169 ( .A(n12095), .ZN(n11969) );
  INV_X1 U9170 ( .A(n8033), .ZN(n6042) );
  INV_X8 U9171 ( .A(n10477), .ZN(n8033) );
  INV_X2 U9172 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U9173 ( .A1(n12448), .A2(n12449), .ZN(n12372) );
  AOI21_X4 U9174 ( .B1(n6435), .B2(n6040), .A(n10832), .ZN(n10740) );
  NAND2_X4 U9175 ( .A1(n11022), .A2(n11021), .ZN(n10855) );
  NAND2_X4 U9176 ( .A1(n5871), .A2(n10637), .ZN(n10617) );
  XNOR2_X2 U9177 ( .A(n6001), .B(n6056), .ZN(n6045) );
  INV_X4 U9178 ( .A(n6045), .ZN(n10871) );
  INV_X4 U9179 ( .A(n6056), .ZN(n6057) );
  INV_X2 U9180 ( .A(n9788), .ZN(n7969) );
  NAND3_X2 U9181 ( .A1(n11423), .A2(n11424), .A3(n11422), .ZN(n6047) );
  AND3_X2 U9182 ( .A1(n10905), .A2(n11232), .A3(n10723), .ZN(n10687) );
  XNOR2_X2 U9183 ( .A(n6419), .B(n6511), .ZN(n6049) );
  XNOR2_X2 U9184 ( .A(n5992), .B(n6517), .ZN(n6050) );
  INV_X2 U9185 ( .A(n10928), .ZN(n10930) );
  NAND3_X2 U9186 ( .A1(n11334), .A2(n11333), .A3(n11740), .ZN(n11261) );
  INV_X4 U9187 ( .A(n11801), .ZN(n6051) );
  NAND2_X4 U9188 ( .A1(n4998), .A2(n11775), .ZN(n11800) );
  INV_X8 U9189 ( .A(net359459), .ZN(net359451) );
  OAI21_X2 U9190 ( .B1(net361838), .B2(n10806), .A(n5043), .ZN(n10801) );
  INV_X1 U9191 ( .A(n11048), .ZN(n6149) );
  NAND2_X4 U9192 ( .A1(n11447), .A2(n11448), .ZN(n11462) );
  INV_X1 U9193 ( .A(n12532), .ZN(n6053) );
  AND2_X4 U9194 ( .A1(net368781), .A2(net367043), .ZN(n6054) );
  INV_X4 U9195 ( .A(n6054), .ZN(n8085) );
  NAND2_X2 U9196 ( .A1(n11324), .A2(n11547), .ZN(n11343) );
  AOI21_X2 U9197 ( .B1(n12533), .B2(net359481), .A(n12532), .ZN(net359472) );
  NOR2_X2 U9198 ( .A1(n10646), .A2(n10648), .ZN(n10600) );
  XNOR2_X2 U9199 ( .A(n11293), .B(n6526), .ZN(n6058) );
  CLKBUF_X3 U9200 ( .A(n12121), .Z(n6059) );
  NAND2_X4 U9201 ( .A1(n11730), .A2(n5992), .ZN(n11833) );
  OAI211_X2 U9202 ( .C1(n11634), .C2(n11633), .A(n11632), .B(n11631), .ZN(
        n11635) );
  NAND3_X2 U9203 ( .A1(n11618), .A2(n11617), .A3(n11639), .ZN(n11632) );
  NAND4_X2 U9204 ( .A1(net365030), .A2(net365031), .A3(net365032), .A4(
        net365033), .ZN(n10521) );
  AOI21_X4 U9205 ( .B1(n7993), .B2(n8025), .A(n7992), .ZN(net365031) );
  OAI21_X4 U9206 ( .B1(n10983), .B2(n10984), .A(n10982), .ZN(n6061) );
  OAI21_X2 U9207 ( .B1(n10983), .B2(n10984), .A(n10982), .ZN(n11048) );
  AOI21_X4 U9208 ( .B1(n10981), .B2(n11036), .A(n11045), .ZN(n10982) );
  NAND2_X4 U9209 ( .A1(n11372), .A2(n5977), .ZN(n11374) );
  NAND4_X4 U9210 ( .A1(n7564), .A2(n7563), .A3(n7562), .A4(n7561), .ZN(n9832)
         );
  INV_X16 U9211 ( .A(n6544), .ZN(n6545) );
  INV_X2 U9212 ( .A(n6545), .ZN(n10346) );
  NAND2_X4 U9213 ( .A1(n10861), .A2(n10863), .ZN(n10766) );
  INV_X4 U9214 ( .A(n6062), .ZN(n6063) );
  NOR2_X2 U9215 ( .A1(n11676), .A2(n11686), .ZN(n11677) );
  XNOR2_X2 U9216 ( .A(n11426), .B(n11314), .ZN(n6064) );
  INV_X8 U9217 ( .A(n6064), .ZN(n11745) );
  INV_X16 U9218 ( .A(net369206), .ZN(net377464) );
  INV_X1 U9219 ( .A(net375993), .ZN(net377453) );
  INV_X2 U9220 ( .A(net377453), .ZN(net377454) );
  XNOR2_X2 U9221 ( .A(n12537), .B(n12536), .ZN(net377452) );
  NAND2_X4 U9222 ( .A1(n12502), .A2(n11670), .ZN(n11671) );
  NAND2_X4 U9223 ( .A1(n11321), .A2(n11354), .ZN(n11164) );
  INV_X4 U9224 ( .A(n11354), .ZN(n11356) );
  NAND2_X4 U9225 ( .A1(n11166), .A2(n5047), .ZN(n11354) );
  NAND2_X4 U9226 ( .A1(n12087), .A2(n12033), .ZN(n12090) );
  OR3_X2 U9227 ( .A1(n9881), .A2(n9883), .A3(n5960), .ZN(n6066) );
  NOR2_X4 U9228 ( .A1(n10903), .A2(n10912), .ZN(n6067) );
  NAND2_X4 U9229 ( .A1(n11459), .A2(n11460), .ZN(n11550) );
  XNOR2_X2 U9230 ( .A(n12009), .B(n12105), .ZN(n6068) );
  NAND2_X1 U9231 ( .A1(n6060), .A2(n11619), .ZN(n11631) );
  XNOR2_X1 U9232 ( .A(n10967), .B(n10966), .ZN(net377443) );
  XNOR2_X2 U9233 ( .A(n10967), .B(n10966), .ZN(net377444) );
  NAND2_X4 U9234 ( .A1(n10963), .A2(n10962), .ZN(n10967) );
  AOI21_X2 U9235 ( .B1(n6276), .B2(n12380), .A(n12379), .ZN(n12389) );
  BUF_X32 U9236 ( .A(n11669), .Z(n6069) );
  NAND2_X2 U9237 ( .A1(n11327), .A2(net361073), .ZN(n11328) );
  XNOR2_X2 U9238 ( .A(n12398), .B(n12384), .ZN(n6070) );
  INV_X8 U9239 ( .A(n6113), .ZN(n12384) );
  INV_X8 U9240 ( .A(n11114), .ZN(n6071) );
  INV_X8 U9241 ( .A(n11155), .ZN(n11114) );
  NAND3_X2 U9242 ( .A1(net361523), .A2(net361524), .A3(net361437), .ZN(n11155)
         );
  BUF_X8 U9243 ( .A(n8715), .Z(n6072) );
  INV_X4 U9244 ( .A(n6073), .ZN(n6074) );
  NOR3_X4 U9245 ( .A1(n10936), .A2(n6014), .A3(n10935), .ZN(n10944) );
  XNOR2_X2 U9246 ( .A(n11529), .B(n6519), .ZN(n6076) );
  INV_X4 U9247 ( .A(n11623), .ZN(n11625) );
  OAI211_X1 U9248 ( .C1(n12502), .C2(net359550), .A(n12501), .B(net100619), 
        .ZN(n12503) );
  INV_X2 U9249 ( .A(n12503), .ZN(aluBoi_multBoi_N52) );
  INV_X1 U9250 ( .A(n11167), .ZN(n6077) );
  INV_X2 U9251 ( .A(n6077), .ZN(n6078) );
  NAND3_X4 U9252 ( .A1(n11134), .A2(net361372), .A3(n11135), .ZN(n11139) );
  INV_X4 U9253 ( .A(n6134), .ZN(n6080) );
  OAI22_X4 U9254 ( .A1(n11379), .A2(net368462), .B1(n11453), .B2(net368195), 
        .ZN(n6081) );
  XNOR2_X2 U9255 ( .A(n11450), .B(n6092), .ZN(n6082) );
  XNOR2_X2 U9256 ( .A(n11483), .B(n6523), .ZN(n6083) );
  AND3_X2 U9257 ( .A1(net360651), .A2(n5986), .A3(net360620), .ZN(n6084) );
  AOI22_X4 U9258 ( .A1(n6086), .A2(n6087), .B1(n6087), .B2(n11898), .ZN(n6085)
         );
  INV_X4 U9259 ( .A(n11663), .ZN(n6087) );
  AOI22_X4 U9260 ( .A1(n11763), .A2(n11841), .B1(n11838), .B2(n11837), .ZN(
        n11795) );
  XNOR2_X2 U9261 ( .A(n11085), .B(n11086), .ZN(net377373) );
  INV_X4 U9262 ( .A(n10873), .ZN(n6088) );
  INV_X4 U9263 ( .A(n6088), .ZN(n6089) );
  AND2_X4 U9264 ( .A1(net375867), .A2(net367035), .ZN(net365399) );
  XNOR2_X2 U9265 ( .A(n12480), .B(n12559), .ZN(n6090) );
  INV_X8 U9266 ( .A(n6091), .ZN(n6092) );
  NAND2_X4 U9267 ( .A1(n10607), .A2(net361801), .ZN(n6093) );
  NAND2_X4 U9268 ( .A1(n12416), .A2(n6028), .ZN(net359450) );
  XOR2_X2 U9269 ( .A(n11079), .B(n11204), .Z(n6094) );
  OAI22_X4 U9270 ( .A1(n11041), .A2(net368442), .B1(n11331), .B2(net368187), 
        .ZN(n11204) );
  NAND2_X4 U9271 ( .A1(n11218), .A2(n11219), .ZN(n11226) );
  XNOR2_X2 U9272 ( .A(n11384), .B(n11383), .ZN(n6095) );
  INV_X8 U9273 ( .A(n6081), .ZN(n11384) );
  OAI21_X2 U9274 ( .B1(n12325), .B2(net369197), .A(net359788), .ZN(net359555)
         );
  NAND3_X2 U9275 ( .A1(n12433), .A2(n12435), .A3(n12199), .ZN(n12018) );
  OAI22_X2 U9276 ( .A1(n11764), .A2(net368462), .B1(n6050), .B2(net368195), 
        .ZN(n11814) );
  INV_X32 U9277 ( .A(net369232), .ZN(net377337) );
  INV_X32 U9278 ( .A(net369232), .ZN(net377338) );
  XNOR2_X2 U9279 ( .A(n11514), .B(n6099), .ZN(n6098) );
  INV_X4 U9280 ( .A(n6098), .ZN(n11919) );
  XOR2_X1 U9281 ( .A(n11687), .B(n6092), .Z(n6099) );
  AOI21_X2 U9282 ( .B1(n5553), .B2(n7560), .A(net365399), .ZN(n7561) );
  XNOR2_X2 U9283 ( .A(n11257), .B(n6101), .ZN(n6100) );
  XOR2_X2 U9284 ( .A(n6119), .B(n11274), .Z(n6101) );
  AOI21_X4 U9285 ( .B1(n11815), .B2(n11783), .A(n11821), .ZN(n11781) );
  AOI22_X2 U9286 ( .A1(net368466), .A2(n6535), .B1(n10891), .B2(n10895), .ZN(
        n10902) );
  INV_X1 U9287 ( .A(n6535), .ZN(n10998) );
  INV_X4 U9288 ( .A(net367009), .ZN(net366997) );
  INV_X16 U9289 ( .A(net366995), .ZN(net366965) );
  NAND2_X1 U9290 ( .A1(net359535), .A2(net360273), .ZN(net360279) );
  NOR2_X2 U9291 ( .A1(n11356), .A2(n11355), .ZN(n11359) );
  NAND2_X2 U9292 ( .A1(n11250), .A2(n6527), .ZN(n6104) );
  NAND2_X4 U9293 ( .A1(n6102), .A2(n6103), .ZN(n6105) );
  NAND2_X4 U9294 ( .A1(n6104), .A2(n6105), .ZN(n11295) );
  INV_X4 U9295 ( .A(n11250), .ZN(n6102) );
  INV_X1 U9296 ( .A(n6527), .ZN(n6103) );
  INV_X1 U9297 ( .A(n5204), .ZN(n6106) );
  AOI21_X2 U9298 ( .B1(n12316), .B2(n12315), .A(n10669), .ZN(n10677) );
  AOI21_X2 U9299 ( .B1(n10671), .B2(n10667), .A(n10651), .ZN(n10673) );
  NAND2_X1 U9300 ( .A1(regBoiz_regfile_17__28_), .A2(n6706), .ZN(n853) );
  NOR3_X2 U9301 ( .A1(n6042), .A2(n10475), .A3(n10476), .ZN(n10481) );
  NAND2_X2 U9302 ( .A1(n10605), .A2(n6543), .ZN(n10614) );
  NAND2_X2 U9303 ( .A1(n7670), .A2(n7556), .ZN(n6109) );
  NOR2_X4 U9304 ( .A1(n12029), .A2(n12100), .ZN(n12037) );
  NOR2_X1 U9305 ( .A1(ifInst[0]), .A2(n13343), .ZN(n13345) );
  OAI21_X1 U9306 ( .B1(ifInst[1]), .B2(ifInst[0]), .A(n6581), .ZN(n13339) );
  NOR2_X1 U9307 ( .A1(ifInst[5]), .A2(ifInst[0]), .ZN(n13503) );
  NAND2_X1 U9308 ( .A1(ifInst[0]), .A2(ifInst[1]), .ZN(n13367) );
  NAND4_X1 U9309 ( .A1(ifOut_95_), .A2(ifOut_94_), .A3(n9938), .A4(n9939), 
        .ZN(n9947) );
  AOI21_X1 U9310 ( .B1(n5557), .B2(n9939), .A(ifOut_95_), .ZN(n9944) );
  NAND2_X1 U9311 ( .A1(ifInst[0]), .A2(n6582), .ZN(n13414) );
  XNOR2_X1 U9312 ( .A(n10349), .B(n10348), .ZN(n10354) );
  XNOR2_X1 U9313 ( .A(n10168), .B(n5737), .ZN(n10169) );
  XNOR2_X1 U9314 ( .A(n10194), .B(n5738), .ZN(n10195) );
  XOR2_X1 U9315 ( .A(ifOut_64_), .B(ifInst[0]), .Z(n10407) );
  INV_X8 U9316 ( .A(n9939), .ZN(n10001) );
  NAND2_X1 U9317 ( .A1(ifInst[0]), .A2(n13499), .ZN(n13302) );
  NAND2_X4 U9318 ( .A1(ifOut_64_), .A2(idBoi_temPC_0_), .ZN(n10397) );
  NAND3_X2 U9319 ( .A1(net360651), .A2(n5986), .A3(net360620), .ZN(n11683) );
  NOR2_X1 U9320 ( .A1(n10841), .A2(n10618), .ZN(n10620) );
  INV_X1 U9321 ( .A(n10841), .ZN(n10621) );
  INV_X8 U9322 ( .A(n11163), .ZN(n11319) );
  NAND2_X1 U9323 ( .A1(regBoiz_regfile_22__5_), .A2(net376076), .ZN(n6111) );
  NAND2_X1 U9324 ( .A1(regBoiz_regfile_30__5_), .A2(net376063), .ZN(n6112) );
  NAND2_X2 U9325 ( .A1(n6111), .A2(n6112), .ZN(n7130) );
  MUX2_X2 U9326 ( .A(n7131), .B(n7130), .S(net366967), .Z(n7132) );
  NAND2_X4 U9327 ( .A1(n6085), .A2(n11835), .ZN(n12120) );
  NAND3_X2 U9328 ( .A1(n7766), .A2(n7765), .A3(n7764), .ZN(n7768) );
  NOR3_X1 U9329 ( .A1(n5449), .A2(n7742), .A3(net368548), .ZN(n7769) );
  INV_X1 U9330 ( .A(net368584), .ZN(net360445) );
  NAND2_X4 U9331 ( .A1(n6185), .A2(n11417), .ZN(n11410) );
  NAND3_X2 U9332 ( .A1(n12105), .A2(n12104), .A3(n12024), .ZN(n12244) );
  NAND2_X2 U9333 ( .A1(n12103), .A2(n12104), .ZN(n12106) );
  INV_X8 U9334 ( .A(n5903), .ZN(n6113) );
  NOR2_X2 U9335 ( .A1(net377531), .A2(net360821), .ZN(n6114) );
  INV_X4 U9336 ( .A(n6114), .ZN(n6115) );
  AND2_X2 U9337 ( .A1(n10547), .A2(net362159), .ZN(n6116) );
  NOR2_X4 U9338 ( .A1(n6116), .A2(net362216), .ZN(net362061) );
  NAND2_X2 U9339 ( .A1(n10518), .A2(net361801), .ZN(n10519) );
  OAI21_X1 U9340 ( .B1(net362211), .B2(n10546), .A(n10545), .ZN(n10547) );
  INV_X1 U9341 ( .A(n10455), .ZN(n6117) );
  INV_X8 U9342 ( .A(n12449), .ZN(n12385) );
  OAI21_X1 U9343 ( .B1(net368181), .B2(n11833), .A(n11832), .ZN(n12096) );
  NAND2_X1 U9344 ( .A1(regBoiz_regfile_27__18_), .A2(n6745), .ZN(n496) );
  NAND2_X2 U9345 ( .A1(n6423), .A2(n11273), .ZN(n6120) );
  NAND2_X4 U9346 ( .A1(n6118), .A2(n6119), .ZN(n6121) );
  NAND2_X4 U9347 ( .A1(n6121), .A2(n6120), .ZN(n11275) );
  INV_X4 U9348 ( .A(n11273), .ZN(n6118) );
  INV_X2 U9349 ( .A(n4988), .ZN(n6122) );
  NAND2_X4 U9350 ( .A1(n10631), .A2(n10688), .ZN(n10632) );
  OAI21_X2 U9351 ( .B1(n11765), .B2(n6517), .A(net368584), .ZN(n11774) );
  NAND3_X2 U9352 ( .A1(n11365), .A2(n11352), .A3(n4996), .ZN(net361021) );
  NAND2_X1 U9353 ( .A1(n10658), .A2(n10657), .ZN(n10660) );
  NAND2_X4 U9354 ( .A1(n7956), .A2(n9867), .ZN(n7961) );
  NAND2_X4 U9355 ( .A1(n11218), .A2(n11219), .ZN(n11222) );
  INV_X32 U9356 ( .A(n6792), .ZN(n6787) );
  INV_X32 U9357 ( .A(n6797), .ZN(n6790) );
  XNOR2_X1 U9358 ( .A(n9106), .B(n6052), .ZN(n13029) );
  AOI21_X1 U9359 ( .B1(n9106), .B2(n6052), .A(n9104), .ZN(n9107) );
  OAI21_X1 U9360 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9071) );
  AOI21_X1 U9361 ( .B1(n9096), .B2(n9095), .A(n9094), .ZN(n9099) );
  INV_X1 U9362 ( .A(n8875), .ZN(n8878) );
  NOR2_X1 U9363 ( .A1(n12094), .A2(n12095), .ZN(n12097) );
  INV_X1 U9364 ( .A(net368584), .ZN(net360205) );
  NAND2_X2 U9365 ( .A1(n12085), .A2(n12418), .ZN(n12137) );
  INV_X32 U9366 ( .A(net366905), .ZN(net377166) );
  INV_X2 U9367 ( .A(n12368), .ZN(n6123) );
  INV_X1 U9368 ( .A(n12275), .ZN(n6124) );
  INV_X2 U9369 ( .A(n6436), .ZN(n6437) );
  NAND2_X1 U9370 ( .A1(regBoiz_regfile_4__29_), .A2(net376417), .ZN(n6125) );
  NAND2_X2 U9371 ( .A1(n6125), .A2(n6126), .ZN(net364970) );
  INV_X4 U9372 ( .A(net368501), .ZN(net368502) );
  XOR2_X1 U9373 ( .A(n6089), .B(n10874), .Z(n10867) );
  NAND2_X2 U9374 ( .A1(n10585), .A2(n10587), .ZN(net376960) );
  INV_X4 U9375 ( .A(n10651), .ZN(n6127) );
  INV_X2 U9376 ( .A(n10650), .ZN(n10651) );
  OAI211_X4 U9377 ( .C1(net361076), .C2(net361077), .A(n5985), .B(n11367), 
        .ZN(n11357) );
  NOR2_X4 U9378 ( .A1(n11512), .A2(n11513), .ZN(n6128) );
  INV_X4 U9379 ( .A(n6128), .ZN(n11509) );
  INV_X4 U9380 ( .A(n11648), .ZN(n6129) );
  NAND2_X4 U9381 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  INV_X4 U9382 ( .A(n10535), .ZN(n6130) );
  NOR2_X2 U9383 ( .A1(n10824), .A2(n10823), .ZN(n10737) );
  BUF_X8 U9384 ( .A(net362230), .Z(net377133) );
  INV_X2 U9385 ( .A(n10544), .ZN(n10546) );
  XNOR2_X1 U9386 ( .A(n9735), .B(n9736), .ZN(n9739) );
  INV_X4 U9387 ( .A(n12479), .ZN(n12559) );
  NAND2_X2 U9388 ( .A1(n12418), .A2(n12153), .ZN(n6131) );
  NAND2_X4 U9389 ( .A1(n12419), .A2(n6132), .ZN(n12375) );
  INV_X4 U9390 ( .A(n6131), .ZN(n6132) );
  NOR2_X2 U9391 ( .A1(n10475), .A2(n10476), .ZN(n8034) );
  INV_X16 U9392 ( .A(n6797), .ZN(n6792) );
  INV_X32 U9393 ( .A(n6798), .ZN(n6797) );
  NAND2_X1 U9394 ( .A1(net368201), .A2(n4999), .ZN(n10904) );
  NAND2_X4 U9395 ( .A1(n8876), .A2(n8875), .ZN(n8879) );
  NAND2_X2 U9396 ( .A1(n6133), .A2(n6134), .ZN(n6136) );
  INV_X1 U9397 ( .A(n10761), .ZN(n6133) );
  NAND2_X4 U9398 ( .A1(n12463), .A2(n12359), .ZN(n12076) );
  NAND2_X4 U9399 ( .A1(n12391), .A2(n12392), .ZN(n12381) );
  NAND2_X1 U9400 ( .A1(regBoiz_regfile_3__28_), .A2(n6492), .ZN(n6137) );
  NAND2_X2 U9401 ( .A1(n6137), .A2(n6138), .ZN(n8000) );
  NAND2_X4 U9402 ( .A1(n8034), .A2(n8033), .ZN(n6147) );
  INV_X4 U9403 ( .A(n6399), .ZN(n6139) );
  INV_X4 U9404 ( .A(n12464), .ZN(n6399) );
  XNOR2_X2 U9405 ( .A(n12241), .B(n12240), .ZN(n12301) );
  AOI21_X4 U9406 ( .B1(net376877), .B2(net362318), .A(net362047), .ZN(
        net362312) );
  INV_X2 U9407 ( .A(n11136), .ZN(n11134) );
  INV_X4 U9408 ( .A(n11033), .ZN(n11129) );
  NOR2_X4 U9409 ( .A1(net360017), .A2(n5558), .ZN(net377071) );
  OAI21_X4 U9410 ( .B1(n7969), .B2(n5872), .A(net362297), .ZN(n10563) );
  AOI22_X4 U9411 ( .A1(n10790), .A2(n10789), .B1(n10792), .B2(net368211), .ZN(
        n10834) );
  NAND2_X4 U9412 ( .A1(n11264), .A2(n5939), .ZN(n11268) );
  NAND2_X4 U9413 ( .A1(n12504), .A2(net378220), .ZN(n11682) );
  NAND2_X4 U9414 ( .A1(n11169), .A2(aluBoi_multBoi_temppp[40]), .ZN(net359923)
         );
  NAND3_X4 U9415 ( .A1(n6392), .A2(n5937), .A3(n12392), .ZN(n12397) );
  INV_X8 U9416 ( .A(n11682), .ZN(n12330) );
  NAND3_X2 U9417 ( .A1(n5933), .A2(n11663), .A3(n11662), .ZN(n11835) );
  MUX2_X2 U9418 ( .A(n6141), .B(n6142), .S(net375867), .Z(n6140) );
  INV_X2 U9419 ( .A(net362270), .ZN(net362269) );
  XNOR2_X2 U9420 ( .A(n12367), .B(n5041), .ZN(n6143) );
  XNOR2_X2 U9421 ( .A(n12145), .B(n12146), .ZN(net359681) );
  NAND2_X2 U9422 ( .A1(n12368), .A2(n12393), .ZN(n12247) );
  INV_X4 U9423 ( .A(n12247), .ZN(n12422) );
  INV_X8 U9424 ( .A(n11707), .ZN(n11389) );
  INV_X8 U9425 ( .A(n10696), .ZN(n10905) );
  AOI21_X2 U9426 ( .B1(n12562), .B2(n12563), .A(n12561), .ZN(n12564) );
  INV_X2 U9427 ( .A(n11268), .ZN(n11266) );
  NAND2_X4 U9428 ( .A1(n11509), .A2(n11508), .ZN(n11515) );
  OAI22_X2 U9429 ( .A1(net362153), .A2(net362134), .B1(n6130), .B2(n10583), 
        .ZN(n10584) );
  NAND2_X1 U9430 ( .A1(n11571), .A2(n11544), .ZN(n6152) );
  NAND2_X4 U9431 ( .A1(n10572), .A2(n10616), .ZN(n10634) );
  NAND2_X4 U9432 ( .A1(n10576), .A2(n10616), .ZN(n10635) );
  NAND2_X2 U9433 ( .A1(n10573), .A2(n6543), .ZN(n10574) );
  OAI21_X2 U9434 ( .B1(n5683), .B2(n6775), .A(n109), .ZN(n4497) );
  INV_X4 U9435 ( .A(n12031), .ZN(n12032) );
  INV_X4 U9436 ( .A(n11410), .ZN(n11494) );
  NAND2_X2 U9437 ( .A1(n11598), .A2(n5213), .ZN(n11599) );
  INV_X1 U9438 ( .A(n11224), .ZN(n11215) );
  NAND2_X1 U9439 ( .A1(net359603), .A2(net368584), .ZN(n11974) );
  NAND3_X1 U9440 ( .A1(n12173), .A2(n12172), .A3(n12256), .ZN(n12180) );
  NAND3_X2 U9441 ( .A1(n10939), .A2(n11096), .A3(n6014), .ZN(n10940) );
  OAI21_X4 U9442 ( .B1(n10943), .B2(n10941), .A(n10940), .ZN(n10942) );
  INV_X4 U9443 ( .A(n12014), .ZN(n11845) );
  NAND4_X2 U9444 ( .A1(n10970), .A2(n10952), .A3(n10953), .A4(net361629), .ZN(
        n11035) );
  NAND2_X2 U9445 ( .A1(n10996), .A2(n6067), .ZN(n10999) );
  NOR2_X4 U9446 ( .A1(n12443), .A2(n12442), .ZN(n12445) );
  AOI22_X4 U9447 ( .A1(regBoiz_regfile_12__12_), .A2(net367003), .B1(
        regBoiz_regfile_14__12_), .B2(net366985), .ZN(n7358) );
  AOI211_X4 U9448 ( .C1(n12432), .C2(n12562), .A(n12431), .B(n12430), .ZN(
        n12443) );
  NAND3_X2 U9449 ( .A1(n11278), .A2(n11049), .A3(n10986), .ZN(n10993) );
  INV_X4 U9450 ( .A(n10954), .ZN(n10961) );
  NAND2_X2 U9451 ( .A1(n10829), .A2(n10841), .ZN(n10957) );
  INV_X4 U9452 ( .A(n11601), .ZN(n11460) );
  OAI22_X1 U9453 ( .A1(n11454), .A2(net368436), .B1(net368179), .B2(n11453), 
        .ZN(n11565) );
  OAI22_X1 U9454 ( .A1(n11454), .A2(net368446), .B1(net368187), .B2(n11453), 
        .ZN(n11502) );
  NOR2_X4 U9455 ( .A1(n12539), .A2(n5009), .ZN(n12547) );
  NAND2_X2 U9456 ( .A1(n11564), .A2(n11563), .ZN(n11685) );
  INV_X2 U9457 ( .A(n11505), .ZN(n11507) );
  OAI22_X1 U9458 ( .A1(n11003), .A2(net368436), .B1(n11331), .B2(net368179), 
        .ZN(n11345) );
  NAND2_X2 U9459 ( .A1(n12392), .A2(n12391), .ZN(n6276) );
  NAND2_X4 U9460 ( .A1(n11579), .A2(n11580), .ZN(n11581) );
  NAND2_X4 U9461 ( .A1(n6145), .A2(n6146), .ZN(net376961) );
  NAND2_X4 U9462 ( .A1(net376960), .A2(net376961), .ZN(n10748) );
  INV_X4 U9463 ( .A(n10585), .ZN(n6145) );
  INV_X1 U9464 ( .A(n10587), .ZN(n6146) );
  NAND3_X2 U9465 ( .A1(n10699), .A2(n11000), .A3(n10698), .ZN(n10700) );
  INV_X2 U9466 ( .A(net359762), .ZN(net359771) );
  INV_X1 U9467 ( .A(n5873), .ZN(n11256) );
  NOR2_X2 U9468 ( .A1(n12119), .A2(n12118), .ZN(n12125) );
  NOR2_X2 U9469 ( .A1(n12468), .A2(n12437), .ZN(n12470) );
  INV_X1 U9470 ( .A(n12557), .ZN(n12560) );
  OAI21_X1 U9471 ( .B1(n6050), .B2(net368181), .A(n12019), .ZN(n12114) );
  OAI22_X1 U9472 ( .A1(n10089), .A2(net368442), .B1(n4992), .B2(net368187), 
        .ZN(n11986) );
  INV_X1 U9473 ( .A(n11785), .ZN(n11787) );
  XNOR2_X2 U9474 ( .A(n11889), .B(n6430), .ZN(n11891) );
  NAND2_X2 U9475 ( .A1(n10582), .A2(net375794), .ZN(n10619) );
  INV_X8 U9476 ( .A(net362152), .ZN(net362196) );
  NOR3_X4 U9477 ( .A1(net366965), .A2(n8123), .A3(n8122), .ZN(n8124) );
  OAI21_X2 U9478 ( .B1(n6624), .B2(n6711), .A(n786), .ZN(n4409) );
  OAI22_X4 U9479 ( .A1(n8051), .A2(net366987), .B1(n8050), .B2(net367003), 
        .ZN(n10446) );
  NOR2_X1 U9480 ( .A1(net360497), .A2(n6573), .ZN(n10080) );
  OAI21_X1 U9481 ( .B1(n6562), .B2(n9525), .A(net368584), .ZN(n9529) );
  OAI21_X1 U9482 ( .B1(net368584), .B2(n6564), .A(n6561), .ZN(n9526) );
  XNOR2_X1 U9483 ( .A(n6113), .B(net359418), .ZN(n12402) );
  NAND2_X1 U9484 ( .A1(n9451), .A2(net368584), .ZN(n9453) );
  XNOR2_X1 U9485 ( .A(net360497), .B(n9451), .ZN(n9736) );
  INV_X16 U9486 ( .A(net368584), .ZN(net360497) );
  NAND2_X4 U9487 ( .A1(net376914), .A2(aluBoi_multBoi_temppp[57]), .ZN(n6148)
         );
  NAND2_X4 U9488 ( .A1(net376916), .A2(n6148), .ZN(net359487) );
  INV_X4 U9489 ( .A(net360033), .ZN(net376914) );
  INV_X4 U9490 ( .A(n6149), .ZN(n6150) );
  NAND2_X4 U9491 ( .A1(n6152), .A2(n6153), .ZN(n11659) );
  NAND2_X4 U9492 ( .A1(n6154), .A2(n6155), .ZN(n6157) );
  NAND2_X4 U9493 ( .A1(n6156), .A2(n6157), .ZN(n12290) );
  INV_X2 U9494 ( .A(n12096), .ZN(n6155) );
  XNOR2_X2 U9495 ( .A(n12290), .B(n5572), .ZN(n12146) );
  NAND2_X2 U9496 ( .A1(n12290), .A2(n12289), .ZN(n12297) );
  NAND4_X4 U9497 ( .A1(n11320), .A2(n11367), .A3(net361088), .A4(n11338), .ZN(
        n11358) );
  NAND2_X2 U9498 ( .A1(n10636), .A2(n10637), .ZN(n10638) );
  NAND3_X2 U9499 ( .A1(n11236), .A2(n11237), .A3(n11235), .ZN(n11310) );
  NOR2_X2 U9500 ( .A1(n6420), .A2(n11607), .ZN(n11521) );
  NAND2_X2 U9501 ( .A1(n12548), .A2(n12551), .ZN(n12487) );
  AOI21_X4 U9502 ( .B1(n12465), .B2(n6139), .A(n5926), .ZN(n12467) );
  OAI21_X4 U9503 ( .B1(n11582), .B2(n11581), .A(n11614), .ZN(n11583) );
  NAND2_X4 U9504 ( .A1(n11884), .A2(n11885), .ZN(n11929) );
  NAND2_X4 U9505 ( .A1(n9089), .A2(n9088), .ZN(n8718) );
  INV_X1 U9506 ( .A(net377133), .ZN(net376877) );
  NAND2_X1 U9507 ( .A1(n11037), .A2(net361443), .ZN(n6160) );
  NAND2_X2 U9508 ( .A1(n6159), .A2(net376879), .ZN(n6161) );
  NAND2_X4 U9509 ( .A1(n6160), .A2(n6161), .ZN(n11125) );
  INV_X2 U9510 ( .A(n11037), .ZN(n6159) );
  INV_X1 U9511 ( .A(net361443), .ZN(net376879) );
  NAND2_X2 U9512 ( .A1(n11912), .A2(n11686), .ZN(n6162) );
  NAND2_X4 U9513 ( .A1(n6163), .A2(n11683), .ZN(net360605) );
  INV_X4 U9514 ( .A(n6162), .ZN(n6163) );
  XNOR2_X2 U9515 ( .A(net377800), .B(net359914), .ZN(n12224) );
  NAND3_X4 U9516 ( .A1(net361808), .A2(net368213), .A3(n10950), .ZN(n10786) );
  OAI21_X4 U9517 ( .B1(n11713), .B2(n11712), .A(n11711), .ZN(n11715) );
  INV_X4 U9518 ( .A(n11699), .ZN(n11706) );
  OAI21_X2 U9519 ( .B1(n11669), .B2(n5335), .A(net359916), .ZN(n11673) );
  INV_X16 U9520 ( .A(n13530), .ZN(n6536) );
  OAI21_X4 U9521 ( .B1(net368225), .B2(n5491), .A(n7639), .ZN(n13530) );
  OAI21_X4 U9522 ( .B1(n11644), .B2(n11468), .A(n11640), .ZN(n11469) );
  NAND2_X4 U9523 ( .A1(n11413), .A2(n11415), .ZN(n11424) );
  INV_X1 U9524 ( .A(n11494), .ZN(n6164) );
  NAND2_X4 U9525 ( .A1(n10709), .A2(n11229), .ZN(n10710) );
  NOR3_X2 U9526 ( .A1(net368502), .A2(net377531), .A3(net375435), .ZN(n10709)
         );
  INV_X8 U9527 ( .A(n11119), .ZN(n11323) );
  INV_X4 U9528 ( .A(n6188), .ZN(n7779) );
  INV_X4 U9529 ( .A(net362097), .ZN(net362094) );
  NAND2_X4 U9530 ( .A1(n11276), .A2(n5973), .ZN(n11432) );
  INV_X8 U9531 ( .A(n11854), .ZN(n11660) );
  NAND2_X2 U9532 ( .A1(n7781), .A2(n6221), .ZN(n6165) );
  NAND2_X2 U9533 ( .A1(n7780), .A2(n6788), .ZN(n6166) );
  NAND2_X4 U9534 ( .A1(n6186), .A2(n6187), .ZN(n7780) );
  INV_X2 U9535 ( .A(n7803), .ZN(n7806) );
  NAND2_X2 U9536 ( .A1(n11420), .A2(n6100), .ZN(n11490) );
  INV_X2 U9537 ( .A(n10868), .ZN(n10679) );
  NAND2_X1 U9538 ( .A1(n8700), .A2(net362253), .ZN(n13525) );
  NAND2_X4 U9539 ( .A1(n11553), .A2(n11534), .ZN(n11586) );
  NAND2_X1 U9540 ( .A1(n10586), .A2(n6093), .ZN(net362124) );
  INV_X2 U9541 ( .A(n10586), .ZN(n10469) );
  AOI21_X2 U9542 ( .B1(net359521), .B2(n12517), .A(n12516), .ZN(
        aluBoi_multBoi_N60) );
  INV_X2 U9543 ( .A(n11907), .ZN(n11910) );
  NAND2_X2 U9544 ( .A1(n11602), .A2(n6277), .ZN(n11603) );
  INV_X1 U9545 ( .A(n10557), .ZN(n10516) );
  NAND2_X4 U9546 ( .A1(n10939), .A2(n10947), .ZN(n10943) );
  XNOR2_X1 U9547 ( .A(n9044), .B(n9045), .ZN(n13129) );
  MUX2_X2 U9548 ( .A(regBoiz_regfile_14__10_), .B(regBoiz_regfile_15__10_), 
        .S(net369244), .Z(n9018) );
  NAND2_X4 U9549 ( .A1(n6169), .A2(n6170), .ZN(n10841) );
  NAND4_X4 U9550 ( .A1(n10749), .A2(net361903), .A3(net361907), .A4(n10750), 
        .ZN(net361886) );
  NAND2_X1 U9551 ( .A1(n9620), .A2(net377611), .ZN(n9624) );
  NAND2_X1 U9552 ( .A1(net361053), .A2(net361088), .ZN(n11115) );
  AOI21_X2 U9553 ( .B1(n7628), .B2(n7627), .A(net366967), .ZN(n7631) );
  INV_X4 U9554 ( .A(n6798), .ZN(n6796) );
  NAND2_X4 U9555 ( .A1(n11537), .A2(n11536), .ZN(n11614) );
  XNOR2_X2 U9556 ( .A(n11480), .B(n6519), .ZN(n11482) );
  NAND3_X2 U9557 ( .A1(n11479), .A2(n11609), .A3(n11527), .ZN(n11480) );
  OAI211_X4 U9558 ( .C1(n6240), .C2(n6437), .A(n12558), .B(net129670), .ZN(
        net359459) );
  NAND2_X1 U9559 ( .A1(n11118), .A2(n11117), .ZN(n11122) );
  NOR2_X2 U9560 ( .A1(n5963), .A2(n11751), .ZN(n11757) );
  AOI21_X4 U9561 ( .B1(n11554), .B2(n11553), .A(n11552), .ZN(n11555) );
  NOR2_X4 U9562 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  NAND2_X1 U9563 ( .A1(n8768), .A2(n6533), .ZN(n8884) );
  OAI22_X1 U9564 ( .A1(n7356), .A2(net367029), .B1(n7355), .B2(net367043), 
        .ZN(n7360) );
  INV_X8 U9565 ( .A(n11620), .ZN(n11615) );
  AOI22_X2 U9566 ( .A1(regBoiz_regfile_8__12_), .A2(net367003), .B1(
        regBoiz_regfile_10__12_), .B2(net366985), .ZN(n7356) );
  INV_X16 U9567 ( .A(net367007), .ZN(net367003) );
  INV_X4 U9568 ( .A(n10468), .ZN(n10455) );
  INV_X2 U9569 ( .A(n6171), .ZN(n6172) );
  NAND2_X1 U9570 ( .A1(n7211), .A2(net376541), .ZN(n6473) );
  NAND2_X4 U9571 ( .A1(n6007), .A2(net378013), .ZN(net361358) );
  OAI21_X2 U9572 ( .B1(n6266), .B2(n5310), .A(n7031), .ZN(n13707) );
  NAND2_X2 U9573 ( .A1(n6327), .A2(n6328), .ZN(n7308) );
  INV_X8 U9574 ( .A(n6796), .ZN(n6795) );
  NAND3_X4 U9575 ( .A1(n10441), .A2(n10440), .A3(n6782), .ZN(n10442) );
  INV_X8 U9576 ( .A(n11459), .ZN(n11713) );
  NAND2_X2 U9577 ( .A1(n7670), .A2(n7645), .ZN(n7650) );
  INV_X4 U9578 ( .A(n6290), .ZN(n8175) );
  NAND2_X1 U9579 ( .A1(n9877), .A2(n6230), .ZN(n6173) );
  NAND2_X2 U9580 ( .A1(n6173), .A2(n6174), .ZN(n7805) );
  NAND2_X4 U9581 ( .A1(n7796), .A2(n7795), .ZN(n9877) );
  INV_X2 U9582 ( .A(n9469), .ZN(n9472) );
  NAND2_X1 U9583 ( .A1(regBoiz_regfile_30__5_), .A2(n340), .ZN(n345) );
  OAI21_X1 U9584 ( .B1(n12064), .B2(net368185), .A(n11994), .ZN(n12273) );
  NAND2_X4 U9585 ( .A1(n11224), .A2(n11223), .ZN(n11264) );
  NAND2_X1 U9586 ( .A1(regBoiz_regfile_15__23_), .A2(n6699), .ZN(n925) );
  OAI21_X4 U9587 ( .B1(n11265), .B2(n6277), .A(n11400), .ZN(n11078) );
  NOR2_X2 U9588 ( .A1(n9871), .A2(n9870), .ZN(n9872) );
  NOR2_X4 U9589 ( .A1(n6016), .A2(n12415), .ZN(n12411) );
  NAND3_X2 U9590 ( .A1(n11727), .A2(n11726), .A3(n11725), .ZN(n11768) );
  INV_X8 U9591 ( .A(n11469), .ZN(n11553) );
  NAND2_X4 U9592 ( .A1(n5919), .A2(n12014), .ZN(n11885) );
  INV_X4 U9593 ( .A(n10889), .ZN(n9789) );
  OAI21_X1 U9594 ( .B1(n6535), .B2(n6563), .A(n6560), .ZN(n9659) );
  NAND2_X1 U9595 ( .A1(n8450), .A2(n6535), .ZN(n8930) );
  NAND2_X1 U9596 ( .A1(n6535), .A2(n13533), .ZN(n11173) );
  AOI22_X2 U9597 ( .A1(regBoiz_regfile_4__12_), .A2(net367003), .B1(
        regBoiz_regfile_6__12_), .B2(net366985), .ZN(n7352) );
  INV_X2 U9598 ( .A(n6175), .ZN(n6176) );
  NAND2_X1 U9599 ( .A1(regBoiz_regfile_19__28_), .A2(n6712), .ZN(n786) );
  INV_X16 U9600 ( .A(net367039), .ZN(net376222) );
  INV_X16 U9601 ( .A(net367039), .ZN(net367023) );
  NAND2_X2 U9602 ( .A1(n11200), .A2(n11201), .ZN(n6179) );
  NAND2_X4 U9603 ( .A1(n6177), .A2(n6178), .ZN(n6180) );
  NAND2_X4 U9604 ( .A1(n6179), .A2(n6180), .ZN(n11221) );
  INV_X4 U9605 ( .A(n11201), .ZN(n6177) );
  INV_X4 U9606 ( .A(n11200), .ZN(n6178) );
  NAND2_X2 U9607 ( .A1(n11222), .A2(n11225), .ZN(n6183) );
  NAND2_X4 U9608 ( .A1(n6181), .A2(n6182), .ZN(n6184) );
  NAND2_X4 U9609 ( .A1(n6183), .A2(n6184), .ZN(n11373) );
  INV_X4 U9610 ( .A(n11222), .ZN(n6181) );
  INV_X8 U9611 ( .A(n11225), .ZN(n6182) );
  NAND2_X4 U9612 ( .A1(n11221), .A2(n11220), .ZN(n11225) );
  XNOR2_X2 U9613 ( .A(n5246), .B(n11202), .ZN(n6185) );
  OAI21_X2 U9614 ( .B1(n5682), .B2(n6694), .A(n953), .ZN(n4437) );
  NOR2_X4 U9615 ( .A1(n11741), .A2(n11496), .ZN(n11411) );
  OAI21_X2 U9616 ( .B1(n6441), .B2(net375435), .A(n10466), .ZN(n10489) );
  INV_X16 U9617 ( .A(net362337), .ZN(net362256) );
  NAND2_X2 U9618 ( .A1(n7779), .A2(net375547), .ZN(n6186) );
  NAND2_X1 U9619 ( .A1(n7778), .A2(net366973), .ZN(n6187) );
  MUX2_X2 U9620 ( .A(n6189), .B(n6190), .S(regBoiz_N12), .Z(n6188) );
  NAND2_X2 U9621 ( .A1(n7647), .A2(net368862), .ZN(n6191) );
  NAND2_X2 U9622 ( .A1(n7646), .A2(net366971), .ZN(n6192) );
  NAND2_X2 U9623 ( .A1(n6191), .A2(n6192), .ZN(n7648) );
  AOI21_X1 U9624 ( .B1(n5553), .B2(n7648), .A(net365399), .ZN(n7649) );
  INV_X2 U9625 ( .A(net362152), .ZN(net362053) );
  NAND2_X2 U9626 ( .A1(net360904), .A2(n10770), .ZN(n10789) );
  AOI211_X1 U9627 ( .C1(n9676), .C2(n6533), .A(n9675), .B(n9674), .ZN(n13049)
         );
  NAND2_X1 U9628 ( .A1(net359603), .A2(n6533), .ZN(n11262) );
  XNOR2_X1 U9629 ( .A(n8767), .B(n6533), .ZN(n8935) );
  NAND2_X1 U9630 ( .A1(net360821), .A2(n13533), .ZN(n11005) );
  INV_X8 U9631 ( .A(n11296), .ZN(n6193) );
  INV_X16 U9632 ( .A(n6193), .ZN(n6194) );
  NAND3_X2 U9633 ( .A1(n11531), .A2(n11530), .A3(net368213), .ZN(n11447) );
  NAND2_X4 U9634 ( .A1(n6196), .A2(n6197), .ZN(n11365) );
  INV_X1 U9635 ( .A(n11347), .ZN(n6195) );
  INV_X4 U9636 ( .A(n11365), .ZN(n11366) );
  INV_X1 U9637 ( .A(net361801), .ZN(net376579) );
  NAND2_X2 U9638 ( .A1(n12154), .A2(n12155), .ZN(n12081) );
  NAND2_X1 U9639 ( .A1(n11182), .A2(n11180), .ZN(n13527) );
  NOR2_X2 U9640 ( .A1(n6093), .A2(n11301), .ZN(n6198) );
  NAND2_X1 U9641 ( .A1(regBoiz_regfile_21__26_), .A2(net376574), .ZN(n6199) );
  NAND2_X1 U9642 ( .A1(regBoiz_regfile_29__26_), .A2(net369202), .ZN(n6200) );
  NAND2_X2 U9643 ( .A1(n6199), .A2(n6200), .ZN(n7937) );
  NAND2_X2 U9644 ( .A1(n10611), .A2(n10612), .ZN(n6203) );
  NAND2_X4 U9645 ( .A1(n6201), .A2(n6202), .ZN(n6204) );
  NAND2_X4 U9646 ( .A1(n6203), .A2(n6204), .ZN(n10613) );
  INV_X4 U9647 ( .A(n10611), .ZN(n6202) );
  NAND2_X2 U9648 ( .A1(n11849), .A2(n11856), .ZN(n11852) );
  NAND2_X4 U9649 ( .A1(n10760), .A2(n10860), .ZN(n10863) );
  NAND2_X4 U9650 ( .A1(n6271), .A2(n9803), .ZN(n13526) );
  INV_X4 U9651 ( .A(n6270), .ZN(n6271) );
  NAND2_X2 U9652 ( .A1(n10619), .A2(n10588), .ZN(n10585) );
  NAND2_X2 U9653 ( .A1(n11596), .A2(n5232), .ZN(n11600) );
  INV_X8 U9654 ( .A(n11420), .ZN(n11741) );
  OAI21_X1 U9655 ( .B1(n6562), .B2(n9487), .A(n5231), .ZN(n9491) );
  OAI21_X1 U9656 ( .B1(n5231), .B2(n6564), .A(n6561), .ZN(n9488) );
  NAND2_X1 U9657 ( .A1(net359752), .A2(n6519), .ZN(n11585) );
  NAND2_X4 U9658 ( .A1(n10926), .A2(n10925), .ZN(n10927) );
  NOR2_X4 U9659 ( .A1(n11476), .A2(n5899), .ZN(n11291) );
  INV_X4 U9660 ( .A(n10781), .ZN(n9892) );
  NAND2_X1 U9661 ( .A1(regBoiz_regfile_23__29_), .A2(net376541), .ZN(n6205) );
  NAND2_X1 U9662 ( .A1(regBoiz_regfile_31__29_), .A2(net377166), .ZN(n6206) );
  NAND2_X2 U9663 ( .A1(n6205), .A2(n6206), .ZN(n8061) );
  NOR2_X1 U9664 ( .A1(n6782), .A2(n5310), .ZN(n7230) );
  INV_X8 U9665 ( .A(n6143), .ZN(n6240) );
  NAND3_X2 U9666 ( .A1(n11942), .A2(n5925), .A3(aluBoi_multBoi_temppp[53]), 
        .ZN(net360273) );
  NAND2_X2 U9667 ( .A1(n11942), .A2(n5925), .ZN(net360259) );
  INV_X1 U9668 ( .A(n5772), .ZN(n11692) );
  INV_X1 U9669 ( .A(n11703), .ZN(n6207) );
  NOR2_X2 U9670 ( .A1(n12468), .A2(n12469), .ZN(n12438) );
  AOI21_X2 U9671 ( .B1(n11024), .B2(n10855), .A(n5965), .ZN(n11104) );
  AOI22_X1 U9672 ( .A1(n3356), .A2(n6835), .B1(aluRw[4]), .B2(n6609), .ZN(
        n3355) );
  NOR2_X2 U9673 ( .A1(n12429), .A2(n12428), .ZN(n12431) );
  NAND2_X4 U9674 ( .A1(n10782), .A2(n5936), .ZN(n11059) );
  NAND3_X2 U9675 ( .A1(n5050), .A2(n11715), .A3(n11714), .ZN(n6208) );
  NAND3_X2 U9676 ( .A1(n11715), .A2(n11714), .A3(n5050), .ZN(n11754) );
  INV_X8 U9677 ( .A(n10780), .ZN(n10915) );
  NOR2_X2 U9678 ( .A1(n11249), .A2(n10696), .ZN(n10699) );
  NAND2_X4 U9679 ( .A1(n12151), .A2(n12150), .ZN(net359899) );
  INV_X2 U9680 ( .A(n6403), .ZN(n7284) );
  INV_X4 U9681 ( .A(n11889), .ZN(n11903) );
  NAND2_X4 U9682 ( .A1(n11305), .A2(n11187), .ZN(n11188) );
  OAI22_X4 U9683 ( .A1(net360539), .A2(net368462), .B1(n11881), .B2(net368195), 
        .ZN(n11775) );
  INV_X16 U9684 ( .A(net367039), .ZN(net367019) );
  INV_X4 U9685 ( .A(net362317), .ZN(net362230) );
  NAND2_X4 U9686 ( .A1(n5962), .A2(n11171), .ZN(n11089) );
  NAND2_X4 U9687 ( .A1(n11759), .A2(n11758), .ZN(n11838) );
  NAND2_X2 U9688 ( .A1(n8065), .A2(net368862), .ZN(n6209) );
  NAND2_X2 U9689 ( .A1(n8064), .A2(net366977), .ZN(n6210) );
  NAND2_X2 U9690 ( .A1(n6209), .A2(n6210), .ZN(n8066) );
  NAND3_X2 U9691 ( .A1(n10437), .A2(n10436), .A3(net367041), .ZN(n10441) );
  NAND2_X4 U9692 ( .A1(n11978), .A2(n12053), .ZN(n11979) );
  NOR2_X4 U9693 ( .A1(net359447), .A2(net359448), .ZN(n12550) );
  INV_X2 U9694 ( .A(n11368), .ZN(n11369) );
  OAI211_X4 U9695 ( .C1(n6084), .C2(n11695), .A(n11694), .B(n11693), .ZN(
        n11696) );
  INV_X1 U9696 ( .A(n10842), .ZN(n10695) );
  INV_X8 U9697 ( .A(n11249), .ZN(n10610) );
  INV_X8 U9698 ( .A(n10949), .ZN(n10849) );
  NAND3_X2 U9699 ( .A1(n11640), .A2(n11639), .A3(n11638), .ZN(n11651) );
  NAND2_X2 U9700 ( .A1(n11960), .A2(n11959), .ZN(n11954) );
  OAI21_X1 U9701 ( .B1(n11560), .B2(n11577), .A(n11657), .ZN(n11567) );
  NOR2_X2 U9702 ( .A1(n10956), .A2(n10955), .ZN(n10959) );
  NAND2_X4 U9703 ( .A1(n10828), .A2(n10827), .ZN(n10846) );
  INV_X8 U9704 ( .A(n11399), .ZN(n11265) );
  NAND2_X1 U9705 ( .A1(n12403), .A2(n12402), .ZN(n6213) );
  NAND2_X4 U9706 ( .A1(n6211), .A2(n6212), .ZN(n6214) );
  NAND2_X4 U9707 ( .A1(n6213), .A2(n6214), .ZN(net359495) );
  INV_X2 U9708 ( .A(n12403), .ZN(n6211) );
  INV_X2 U9709 ( .A(n11586), .ZN(n11592) );
  NAND2_X1 U9710 ( .A1(n11710), .A2(n11709), .ZN(n11712) );
  NAND2_X2 U9711 ( .A1(n10972), .A2(n6537), .ZN(n10994) );
  AOI21_X2 U9712 ( .B1(net359462), .B2(n6065), .A(net359418), .ZN(n12541) );
  OAI22_X1 U9713 ( .A1(n11812), .A2(net368436), .B1(n5030), .B2(net368179), 
        .ZN(n12157) );
  NOR2_X4 U9714 ( .A1(n11706), .A2(n11840), .ZN(n11763) );
  NAND2_X1 U9715 ( .A1(n11870), .A2(n11871), .ZN(n11873) );
  INV_X2 U9716 ( .A(n6215), .ZN(n6216) );
  NAND2_X2 U9717 ( .A1(n7376), .A2(net376417), .ZN(n6217) );
  NAND2_X1 U9718 ( .A1(n7375), .A2(net368781), .ZN(n6218) );
  NAND2_X2 U9719 ( .A1(n6217), .A2(n6218), .ZN(n7377) );
  INV_X4 U9720 ( .A(n11778), .ZN(n11806) );
  INV_X32 U9721 ( .A(net366901), .ZN(net368781) );
  INV_X8 U9722 ( .A(net367007), .ZN(net367001) );
  NAND3_X2 U9723 ( .A1(n9815), .A2(n9814), .A3(n9813), .ZN(n9816) );
  INV_X8 U9724 ( .A(n9841), .ZN(n11187) );
  NAND2_X4 U9725 ( .A1(n11030), .A2(n10856), .ZN(n10794) );
  NAND2_X1 U9726 ( .A1(regBoiz_regfile_19__24_), .A2(n6788), .ZN(n7819) );
  OAI22_X4 U9727 ( .A1(n7864), .A2(n7863), .B1(n7862), .B2(n7861), .ZN(n9890)
         );
  INV_X16 U9728 ( .A(n13520), .ZN(n6512) );
  NAND2_X4 U9729 ( .A1(n9802), .A2(n9804), .ZN(n13520) );
  OAI22_X4 U9730 ( .A1(n12059), .A2(net368467), .B1(net368211), .B2(n12342), 
        .ZN(n12175) );
  NAND2_X4 U9731 ( .A1(n12058), .A2(n6421), .ZN(n12342) );
  NAND2_X4 U9732 ( .A1(net375650), .A2(n7782), .ZN(n7803) );
  NAND2_X4 U9733 ( .A1(n10571), .A2(n10570), .ZN(n10605) );
  NAND2_X4 U9734 ( .A1(n9798), .A2(n9805), .ZN(net328053) );
  INV_X16 U9735 ( .A(net368583), .ZN(net368584) );
  INV_X16 U9736 ( .A(n13534), .ZN(n6522) );
  NAND2_X4 U9737 ( .A1(n9812), .A2(n9814), .ZN(n13534) );
  INV_X8 U9738 ( .A(n11338), .ZN(n11339) );
  NAND2_X4 U9739 ( .A1(n9965), .A2(n5696), .ZN(n10191) );
  NAND2_X4 U9740 ( .A1(n9980), .A2(n10030), .ZN(n9982) );
  NAND2_X4 U9741 ( .A1(n5017), .A2(n9979), .ZN(n10030) );
  AOI22_X4 U9742 ( .A1(n10255), .A2(n9959), .B1(idOut_98_), .B2(
        aluBoi_imm32w_12_), .ZN(n10243) );
  OAI22_X4 U9743 ( .A1(n6568), .A2(n5505), .B1(n10072), .B2(n10071), .ZN(
        n10061) );
  OAI22_X4 U9744 ( .A1(n6568), .A2(n5504), .B1(n10135), .B2(n10134), .ZN(
        n10128) );
  NAND2_X2 U9745 ( .A1(n7195), .A2(net376387), .ZN(n6219) );
  NAND2_X1 U9746 ( .A1(n7194), .A2(net378321), .ZN(n6220) );
  NAND2_X2 U9747 ( .A1(n6219), .A2(n6220), .ZN(n7196) );
  NAND2_X2 U9748 ( .A1(n7213), .A2(n6221), .ZN(n6222) );
  NAND2_X1 U9749 ( .A1(n7212), .A2(n6789), .ZN(n6223) );
  NAND2_X2 U9750 ( .A1(n6222), .A2(n6223), .ZN(n7214) );
  NAND2_X4 U9751 ( .A1(n11940), .A2(n5975), .ZN(n11943) );
  XNOR2_X2 U9752 ( .A(n11159), .B(net361007), .ZN(net360636) );
  NOR3_X2 U9753 ( .A1(n5265), .A2(net362251), .A3(n5002), .ZN(n10529) );
  NOR2_X4 U9754 ( .A1(n10528), .A2(n10527), .ZN(n10512) );
  NOR3_X4 U9755 ( .A1(n5031), .A2(n5946), .A3(n11721), .ZN(n11728) );
  INV_X4 U9756 ( .A(n11734), .ZN(n11735) );
  INV_X4 U9757 ( .A(n10605), .ZN(n10606) );
  XNOR2_X1 U9758 ( .A(n11736), .B(n11345), .ZN(n11347) );
  INV_X32 U9759 ( .A(net366905), .ZN(net366887) );
  NAND3_X2 U9760 ( .A1(net369287), .A2(n11082), .A3(n11090), .ZN(n11091) );
  NAND2_X4 U9761 ( .A1(n12073), .A2(n12270), .ZN(n12359) );
  NAND2_X4 U9762 ( .A1(n11460), .A2(n11623), .ZN(n11217) );
  NAND2_X2 U9763 ( .A1(n6224), .A2(net361756), .ZN(n6226) );
  INV_X4 U9764 ( .A(n11097), .ZN(n6224) );
  NOR2_X1 U9765 ( .A1(n12288), .A2(n12423), .ZN(n12160) );
  NAND3_X1 U9766 ( .A1(n12002), .A2(n12022), .A3(n12023), .ZN(n12024) );
  NOR2_X4 U9767 ( .A1(n11493), .A2(n11421), .ZN(n11422) );
  NAND2_X1 U9768 ( .A1(regBoiz_regfile_31__12_), .A2(n6757), .ZN(n335) );
  INV_X4 U9769 ( .A(n11429), .ZN(n11513) );
  NAND2_X4 U9770 ( .A1(n11474), .A2(n11468), .ZN(n11642) );
  INV_X8 U9771 ( .A(n11390), .ZN(n11474) );
  NAND2_X4 U9772 ( .A1(n11891), .A2(n11890), .ZN(n12107) );
  NAND2_X4 U9773 ( .A1(n10732), .A2(n10792), .ZN(n10733) );
  NAND3_X4 U9774 ( .A1(net369286), .A2(n11129), .A3(n11113), .ZN(net361398) );
  OAI221_X4 U9775 ( .B1(n12392), .B2(n12376), .C1(n5909), .C2(n12375), .A(
        n12374), .ZN(n12416) );
  INV_X2 U9776 ( .A(net376321), .ZN(net376322) );
  NAND4_X4 U9777 ( .A1(net360620), .A2(n5772), .A3(n11664), .A4(n11675), .ZN(
        n11518) );
  NAND2_X4 U9778 ( .A1(n12074), .A2(n12073), .ZN(n12463) );
  INV_X8 U9779 ( .A(n10913), .ZN(n11244) );
  INV_X8 U9780 ( .A(n11591), .ZN(n11556) );
  NAND2_X4 U9781 ( .A1(n12029), .A2(n12030), .ZN(n12089) );
  NAND2_X4 U9782 ( .A1(n11398), .A2(n11278), .ZN(n11623) );
  OAI21_X2 U9783 ( .B1(n12170), .B2(n12070), .A(n12173), .ZN(n12072) );
  INV_X2 U9784 ( .A(n10897), .ZN(n10891) );
  AOI21_X4 U9785 ( .B1(n5910), .B2(n10764), .A(n10866), .ZN(n10765) );
  INV_X8 U9786 ( .A(n11495), .ZN(n11742) );
  NAND3_X4 U9787 ( .A1(n11138), .A2(n11140), .A3(n11139), .ZN(n11338) );
  NOR2_X2 U9788 ( .A1(n10955), .A2(n5901), .ZN(n10735) );
  NAND2_X4 U9789 ( .A1(n11398), .A2(n11397), .ZN(n11399) );
  NAND2_X1 U9790 ( .A1(regBoiz_regfile_31__29_), .A2(n6757), .ZN(n317) );
  XNOR2_X1 U9791 ( .A(net362311), .B(net362312), .ZN(n10490) );
  MUX2_X1 U9792 ( .A(regBoiz_regfile_11__23_), .B(regBoiz_regfile_15__23_), 
        .S(net366937), .Z(n7776) );
  OAI21_X4 U9793 ( .B1(n11116), .B2(net368195), .A(n10924), .ZN(n10977) );
  NAND2_X4 U9794 ( .A1(n10977), .A2(n10978), .ZN(n10989) );
  XNOR2_X2 U9795 ( .A(n12255), .B(n6229), .ZN(n12063) );
  NAND2_X1 U9796 ( .A1(n11573), .A2(n5928), .ZN(n11489) );
  NAND2_X2 U9797 ( .A1(n11114), .A2(n11125), .ZN(n11128) );
  NAND2_X4 U9798 ( .A1(n6051), .A2(n11786), .ZN(n11777) );
  INV_X4 U9799 ( .A(n11642), .ZN(n11645) );
  NAND2_X4 U9800 ( .A1(net360821), .A2(n13706), .ZN(n10792) );
  NOR3_X2 U9801 ( .A1(n10501), .A2(net362257), .A3(net368209), .ZN(n10503) );
  INV_X16 U9802 ( .A(net367035), .ZN(net375717) );
  NAND2_X2 U9803 ( .A1(n7276), .A2(n6230), .ZN(n6231) );
  NAND2_X1 U9804 ( .A1(n7275), .A2(n6784), .ZN(n6232) );
  NAND2_X2 U9805 ( .A1(n6231), .A2(n6232), .ZN(n7277) );
  INV_X2 U9806 ( .A(n6233), .ZN(n6234) );
  NAND2_X4 U9807 ( .A1(n11720), .A2(n11719), .ZN(net329432) );
  INV_X8 U9808 ( .A(n11608), .ZN(n11718) );
  AND3_X4 U9809 ( .A1(n11479), .A2(n11719), .A3(n11720), .ZN(n11611) );
  NAND2_X2 U9810 ( .A1(n9988), .A2(n9992), .ZN(dpcHold) );
  NAND3_X2 U9811 ( .A1(n7472), .A2(n7471), .A3(n6054), .ZN(n7473) );
  INV_X32 U9812 ( .A(net366945), .ZN(net366925) );
  INV_X4 U9813 ( .A(n9796), .ZN(n11976) );
  NAND2_X2 U9814 ( .A1(n7408), .A2(n6230), .ZN(n6235) );
  NAND2_X1 U9815 ( .A1(n7407), .A2(n6786), .ZN(n6236) );
  NAND2_X2 U9816 ( .A1(n6235), .A2(n6236), .ZN(n7409) );
  INV_X8 U9817 ( .A(n13519), .ZN(n6510) );
  INV_X4 U9818 ( .A(n7060), .ZN(n6274) );
  MUX2_X1 U9819 ( .A(n7055), .B(n7054), .S(net366977), .Z(n7056) );
  INV_X16 U9820 ( .A(net367035), .ZN(net367029) );
  INV_X4 U9821 ( .A(n11992), .ZN(n9901) );
  NAND3_X2 U9822 ( .A1(n11976), .A2(n9900), .A3(n11977), .ZN(n11992) );
  AOI21_X2 U9823 ( .B1(n10286), .B2(n12853), .A(n6434), .ZN(n10319) );
  NAND3_X2 U9824 ( .A1(n9988), .A2(n9992), .A3(n10286), .ZN(n10383) );
  NOR2_X2 U9825 ( .A1(MoLanBoJ), .A2(n9995), .ZN(n10406) );
  INV_X4 U9826 ( .A(n10383), .ZN(n6550) );
  AOI21_X1 U9827 ( .B1(n6571), .B2(n12710), .A(MoLanBoJ), .ZN(n10123) );
  AOI21_X1 U9828 ( .B1(n6571), .B2(n5355), .A(MoLanBoJ), .ZN(n10370) );
  AOI21_X1 U9829 ( .B1(n6571), .B2(n12810), .A(MoLanBoJ), .ZN(n10265) );
  AOI21_X1 U9830 ( .B1(n10286), .B2(n12613), .A(MoLanBoJ), .ZN(n9990) );
  AOI21_X1 U9831 ( .B1(n6571), .B2(n12770), .A(MoLanBoJ), .ZN(n10200) );
  AOI21_X1 U9832 ( .B1(n6571), .B2(n12745), .A(MoLanBoJ), .ZN(n10162) );
  AOI21_X1 U9833 ( .B1(n6571), .B2(n12854), .A(MoLanBoJ), .ZN(n10314) );
  AOI21_X1 U9834 ( .B1(n10286), .B2(n12725), .A(MoLanBoJ), .ZN(n10145) );
  AOI21_X1 U9835 ( .B1(n6571), .B2(n12625), .A(n6434), .ZN(n10011) );
  NAND2_X1 U9836 ( .A1(regBoiz_regfile_31__13_), .A2(n6757), .ZN(n334) );
  INV_X4 U9837 ( .A(net375525), .ZN(net365830) );
  MUX2_X2 U9838 ( .A(n7144), .B(n7145), .S(net375721), .Z(n7146) );
  MUX2_X1 U9839 ( .A(n7147), .B(n7146), .S(net366919), .Z(n7148) );
  INV_X4 U9840 ( .A(n6325), .ZN(n7110) );
  INV_X2 U9841 ( .A(n6480), .ZN(n7109) );
  MUX2_X1 U9842 ( .A(n7110), .B(n7109), .S(net366981), .Z(n7111) );
  INV_X4 U9843 ( .A(n6302), .ZN(n7114) );
  INV_X2 U9844 ( .A(n6489), .ZN(n7113) );
  NAND2_X2 U9845 ( .A1(n7106), .A2(net375614), .ZN(n6237) );
  NAND2_X1 U9846 ( .A1(n7105), .A2(net367029), .ZN(n6238) );
  NAND2_X2 U9847 ( .A1(n6237), .A2(n6238), .ZN(n7120) );
  INV_X4 U9848 ( .A(n6252), .ZN(n7095) );
  INV_X32 U9849 ( .A(net367039), .ZN(net376223) );
  NAND2_X1 U9850 ( .A1(regBoiz_regfile_27__23_), .A2(n6745), .ZN(n490) );
  NAND2_X2 U9851 ( .A1(n7932), .A2(net368862), .ZN(n6241) );
  NAND2_X1 U9852 ( .A1(n7931), .A2(net366973), .ZN(n6242) );
  NOR2_X4 U9853 ( .A1(n11052), .A2(n9822), .ZN(n9825) );
  NAND2_X2 U9854 ( .A1(net362122), .A2(net361913), .ZN(n10591) );
  MUX2_X1 U9855 ( .A(n7406), .B(n7405), .S(net378488), .Z(n7407) );
  INV_X4 U9856 ( .A(n12118), .ZN(n11904) );
  NAND2_X4 U9857 ( .A1(n10776), .A2(n10777), .ZN(n10822) );
  NAND2_X2 U9858 ( .A1(n11034), .A2(n5882), .ZN(n11093) );
  XNOR2_X2 U9859 ( .A(net377576), .B(net362149), .ZN(net362146) );
  NAND2_X4 U9860 ( .A1(n12164), .A2(n12163), .ZN(n12357) );
  XNOR2_X1 U9861 ( .A(n11255), .B(n5873), .ZN(n11315) );
  NAND2_X1 U9862 ( .A1(regBoiz_regfile_29__23_), .A2(n6751), .ZN(n423) );
  INV_X1 U9863 ( .A(n11127), .ZN(n11133) );
  NAND2_X2 U9864 ( .A1(net375713), .A2(n9819), .ZN(n9820) );
  NOR2_X4 U9865 ( .A1(n10524), .A2(n10525), .ZN(n10534) );
  MUX2_X1 U9866 ( .A(n7240), .B(n7239), .S(net366981), .Z(n7241) );
  NAND2_X4 U9867 ( .A1(net368215), .A2(n6535), .ZN(n10894) );
  NAND2_X4 U9868 ( .A1(net368215), .A2(n10894), .ZN(n10897) );
  NAND3_X1 U9869 ( .A1(n7329), .A2(net376541), .A3(net366953), .ZN(n7334) );
  NAND3_X1 U9870 ( .A1(net366937), .A2(n7315), .A3(n5135), .ZN(n7322) );
  NAND2_X1 U9871 ( .A1(regBoiz_regfile_4__23_), .A2(net366907), .ZN(n7784) );
  NAND2_X1 U9872 ( .A1(regBoiz_regfile_6__23_), .A2(net366907), .ZN(n7790) );
  NAND2_X1 U9873 ( .A1(regBoiz_regfile_0__23_), .A2(net366907), .ZN(n7786) );
  NAND2_X1 U9874 ( .A1(regBoiz_regfile_2__23_), .A2(net366907), .ZN(n7792) );
  AOI22_X1 U9875 ( .A1(regBoiz_regfile_2__29_), .A2(net366907), .B1(
        regBoiz_regfile_10__29_), .B2(net368782), .ZN(n8050) );
  OAI21_X1 U9876 ( .B1(net361891), .B2(net361536), .A(net361827), .ZN(n10756)
         );
  AOI21_X4 U9877 ( .B1(n10523), .B2(n10522), .A(net362262), .ZN(n10524) );
  AOI21_X2 U9878 ( .B1(n11123), .B2(net361372), .A(net361390), .ZN(n11140) );
  INV_X4 U9879 ( .A(n6362), .ZN(n7797) );
  INV_X4 U9880 ( .A(n11635), .ZN(n11711) );
  NAND3_X4 U9881 ( .A1(n11445), .A2(n11446), .A3(n11444), .ZN(n11646) );
  NOR2_X2 U9882 ( .A1(n11303), .A2(n11302), .ZN(n11306) );
  NAND3_X2 U9883 ( .A1(n9840), .A2(n9839), .A3(n9838), .ZN(n11302) );
  NAND2_X4 U9884 ( .A1(n10813), .A2(n10812), .ZN(n10884) );
  NAND3_X2 U9885 ( .A1(n10811), .A2(n10849), .A3(n10950), .ZN(n10812) );
  NAND2_X4 U9886 ( .A1(n10886), .A2(n10885), .ZN(n10950) );
  NAND2_X2 U9887 ( .A1(daddr[2]), .A2(net364968), .ZN(n10451) );
  AOI21_X1 U9888 ( .B1(n7786), .B2(n7785), .A(net366927), .ZN(n7787) );
  OAI21_X1 U9889 ( .B1(n6782), .B2(n5597), .A(net366927), .ZN(n8151) );
  OAI21_X1 U9890 ( .B1(n6782), .B2(n5598), .A(net366927), .ZN(n8153) );
  AOI21_X1 U9891 ( .B1(n7869), .B2(n7868), .A(net366927), .ZN(n7870) );
  NAND3_X2 U9892 ( .A1(n12265), .A2(n12264), .A3(n12263), .ZN(n12266) );
  INV_X8 U9893 ( .A(n10450), .ZN(n10457) );
  INV_X2 U9894 ( .A(net361913), .ZN(net361911) );
  NAND2_X4 U9895 ( .A1(n12275), .A2(n12273), .ZN(n12073) );
  NAND2_X4 U9896 ( .A1(n11126), .A2(n11125), .ZN(n11127) );
  NAND2_X4 U9897 ( .A1(n11160), .A2(n11167), .ZN(n11162) );
  NAND2_X1 U9898 ( .A1(n11230), .A2(n11229), .ZN(n11311) );
  INV_X8 U9899 ( .A(net328053), .ZN(net368583) );
  INV_X8 U9900 ( .A(n11843), .ZN(n11548) );
  INV_X1 U9901 ( .A(n10770), .ZN(n10701) );
  OAI21_X4 U9902 ( .B1(n10947), .B2(n11096), .A(n5882), .ZN(n10948) );
  AOI22_X4 U9903 ( .A1(n11137), .A2(n5334), .B1(n11136), .B2(n5334), .ZN(
        n11138) );
  INV_X8 U9904 ( .A(n10629), .ZN(n10838) );
  NAND2_X4 U9905 ( .A1(n11844), .A2(n11879), .ZN(n6244) );
  NAND2_X4 U9906 ( .A1(n12113), .A2(n6048), .ZN(n12030) );
  OAI21_X4 U9907 ( .B1(n11828), .B2(n11827), .A(n11826), .ZN(n12039) );
  NAND2_X4 U9908 ( .A1(n11724), .A2(n5309), .ZN(n11730) );
  OAI211_X4 U9909 ( .C1(n12001), .C2(n12000), .A(n6002), .B(n5042), .ZN(n12023) );
  INV_X2 U9910 ( .A(n11997), .ZN(n12001) );
  NAND3_X2 U9911 ( .A1(n11029), .A2(n11030), .A3(n11028), .ZN(n11024) );
  AOI21_X1 U9912 ( .B1(n11029), .B2(n11030), .A(n11028), .ZN(n11032) );
  NOR2_X2 U9913 ( .A1(net361416), .A2(n11026), .ZN(n11040) );
  NAND2_X4 U9914 ( .A1(n11933), .A2(net360299), .ZN(n12093) );
  INV_X8 U9915 ( .A(n11518), .ZN(n11933) );
  OAI211_X4 U9916 ( .C1(n11919), .C2(n11918), .A(n11917), .B(n11923), .ZN(
        n11927) );
  NAND2_X2 U9917 ( .A1(n10558), .A2(n10559), .ZN(n6247) );
  NAND2_X4 U9918 ( .A1(n6245), .A2(n6246), .ZN(n6248) );
  NAND2_X4 U9919 ( .A1(n6247), .A2(n6248), .ZN(net362152) );
  INV_X4 U9920 ( .A(n10558), .ZN(n6246) );
  XNOR2_X2 U9921 ( .A(n11847), .B(n11848), .ZN(n6249) );
  NAND2_X4 U9922 ( .A1(n11933), .A2(net360299), .ZN(n12031) );
  NAND2_X4 U9923 ( .A1(n10755), .A2(net361893), .ZN(n10861) );
  NAND2_X1 U9924 ( .A1(net376374), .A2(net366987), .ZN(n8152) );
  NOR3_X4 U9925 ( .A1(net361746), .A2(net361748), .A3(net376691), .ZN(n10857)
         );
  AOI21_X4 U9926 ( .B1(n11788), .B2(n11787), .A(n11802), .ZN(n11789) );
  INV_X8 U9927 ( .A(n10560), .ZN(n6250) );
  MUX2_X2 U9928 ( .A(n6253), .B(n6254), .S(net375867), .Z(n6252) );
  INV_X8 U9929 ( .A(n11723), .ZN(n11528) );
  MUX2_X2 U9930 ( .A(n6462), .B(n6256), .S(net376642), .Z(n6255) );
  MUX2_X2 U9931 ( .A(n7178), .B(n7177), .S(net366933), .Z(n7179) );
  NAND2_X2 U9932 ( .A1(n7100), .A2(net368862), .ZN(n6257) );
  NAND2_X1 U9933 ( .A1(net366184), .A2(net366979), .ZN(n6258) );
  NAND2_X2 U9934 ( .A1(n6257), .A2(n6258), .ZN(n7104) );
  MUX2_X1 U9935 ( .A(n7104), .B(n7103), .S(net366939), .Z(n7105) );
  NAND2_X1 U9936 ( .A1(regBoiz_regfile_4__4_), .A2(net376417), .ZN(n6259) );
  NAND2_X1 U9937 ( .A1(n6320), .A2(net376063), .ZN(n6260) );
  NAND2_X2 U9938 ( .A1(n6259), .A2(n6260), .ZN(n7097) );
  MUX2_X1 U9939 ( .A(n7097), .B(n7096), .S(net366979), .Z(n7098) );
  NAND2_X2 U9940 ( .A1(n7164), .A2(net376387), .ZN(n6261) );
  NAND2_X1 U9941 ( .A1(n7163), .A2(net366939), .ZN(n6262) );
  NAND2_X2 U9942 ( .A1(n6261), .A2(n6262), .ZN(n7165) );
  NAND2_X2 U9943 ( .A1(n7176), .A2(net368862), .ZN(n6263) );
  NAND2_X1 U9944 ( .A1(n7175), .A2(net366967), .ZN(n6264) );
  NAND2_X2 U9945 ( .A1(n6263), .A2(n6264), .ZN(n7177) );
  OAI21_X2 U9946 ( .B1(n5684), .B2(n6755), .A(n310), .ZN(n3695) );
  MUX2_X1 U9947 ( .A(regBoiz_regfile_30__6_), .B(regBoiz_regfile_31__6_), .S(
        net367029), .Z(n7175) );
  MUX2_X1 U9948 ( .A(regBoiz_regfile_14__6_), .B(regBoiz_regfile_15__6_), .S(
        net375717), .Z(n7161) );
  INV_X4 U9949 ( .A(n7030), .ZN(n6267) );
  INV_X4 U9950 ( .A(n7029), .ZN(n6268) );
  INV_X8 U9951 ( .A(n6334), .ZN(n6335) );
  INV_X8 U9952 ( .A(net367035), .ZN(net367031) );
  INV_X8 U9953 ( .A(net367035), .ZN(net367025) );
  MUX2_X2 U9954 ( .A(n6267), .B(n6268), .S(n6785), .Z(n6266) );
  NAND2_X1 U9955 ( .A1(regBoiz_regfile_7__1_), .A2(n6774), .ZN(n156) );
  MUX2_X2 U9956 ( .A(regBoiz_regfile_6__1_), .B(regBoiz_regfile_7__1_), .S(
        net369163), .Z(n9211) );
  MUX2_X1 U9957 ( .A(n7004), .B(n7003), .S(net366977), .Z(n7005) );
  OAI21_X2 U9958 ( .B1(n6272), .B2(n5310), .A(n7062), .ZN(n13519) );
  INV_X4 U9959 ( .A(n7061), .ZN(n6273) );
  MUX2_X1 U9960 ( .A(n7006), .B(n7005), .S(net366933), .Z(n7014) );
  INV_X1 U9961 ( .A(n9797), .ZN(n6270) );
  INV_X4 U9962 ( .A(n6301), .ZN(n7115) );
  INV_X16 U9963 ( .A(net367035), .ZN(net375650) );
  MUX2_X2 U9964 ( .A(n6273), .B(n6274), .S(n6784), .Z(n6272) );
  INV_X2 U9965 ( .A(n11836), .ZN(n6275) );
  INV_X8 U9966 ( .A(n10845), .ZN(n10956) );
  INV_X4 U9967 ( .A(n12133), .ZN(n12138) );
  OAI21_X4 U9968 ( .B1(n11442), .B2(n11491), .A(n5976), .ZN(n11450) );
  INV_X8 U9969 ( .A(n11360), .ZN(n12502) );
  INV_X8 U9970 ( .A(n11271), .ZN(n6277) );
  INV_X1 U9971 ( .A(n12353), .ZN(n12345) );
  NAND2_X2 U9972 ( .A1(n11208), .A2(n11209), .ZN(n11210) );
  NAND2_X1 U9973 ( .A1(net360904), .A2(n5873), .ZN(n11220) );
  NAND2_X1 U9974 ( .A1(net360821), .A2(n5873), .ZN(n11065) );
  NAND3_X4 U9975 ( .A1(n11376), .A2(n5034), .A3(n5939), .ZN(n11377) );
  OAI22_X2 U9976 ( .A1(n12251), .A2(net368462), .B1(n5878), .B2(net368195), 
        .ZN(n12253) );
  OAI22_X4 U9977 ( .A1(n12184), .A2(net368467), .B1(n5878), .B2(net368211), 
        .ZN(n12252) );
  OAI21_X4 U9978 ( .B1(n12253), .B2(n4991), .A(n12573), .ZN(n12460) );
  OAI21_X2 U9979 ( .B1(n5878), .B2(net368185), .A(n12343), .ZN(n12473) );
  OAI21_X2 U9980 ( .B1(n5450), .B2(n7470), .A(net366967), .ZN(n7471) );
  XNOR2_X2 U9981 ( .A(net360259), .B(aluBoi_multBoi_temppp[53]), .ZN(net375993) );
  AOI22_X4 U9982 ( .A1(n8084), .A2(n8083), .B1(n8082), .B2(n8081), .ZN(n8086)
         );
  NAND2_X4 U9983 ( .A1(n12501), .A2(net360628), .ZN(n12328) );
  NAND2_X4 U9984 ( .A1(aluBoi_multBoi_temppp[46]), .A2(n11369), .ZN(net360628)
         );
  NAND2_X4 U9985 ( .A1(n8038), .A2(n8037), .ZN(n10479) );
  NAND2_X4 U9986 ( .A1(n10479), .A2(n10478), .ZN(n10527) );
  AOI21_X4 U9987 ( .B1(n12411), .B2(n12410), .A(n12409), .ZN(n12412) );
  NAND3_X4 U9988 ( .A1(n9788), .A2(n9787), .A3(n10562), .ZN(n10567) );
  NAND2_X4 U9989 ( .A1(n11709), .A2(n11389), .ZN(n11601) );
  INV_X1 U9990 ( .A(n10451), .ZN(n10452) );
  AOI21_X2 U9991 ( .B1(n12295), .B2(n12294), .A(n12293), .ZN(n12296) );
  NAND2_X4 U9992 ( .A1(n10768), .A2(n10769), .ZN(n11103) );
  NAND2_X4 U9993 ( .A1(n11029), .A2(n11030), .ZN(n10768) );
  INV_X8 U9994 ( .A(n6194), .ZN(n6279) );
  INV_X4 U9995 ( .A(n6280), .ZN(n7192) );
  MUX2_X2 U9996 ( .A(n7193), .B(n7192), .S(net375527), .Z(n7194) );
  NAND2_X4 U9997 ( .A1(n7944), .A2(net366953), .ZN(n7990) );
  INV_X2 U9998 ( .A(n7990), .ZN(n7934) );
  OAI211_X1 U9999 ( .C1(n6787), .C2(n5590), .A(n8127), .B(net366953), .ZN(
        n8130) );
  NAND2_X4 U10000 ( .A1(n8069), .A2(net366953), .ZN(n10437) );
  MUX2_X2 U10001 ( .A(n6454), .B(n6281), .S(net367043), .Z(n6280) );
  INV_X1 U10002 ( .A(n10552), .ZN(n6282) );
  INV_X2 U10003 ( .A(n6283), .ZN(n6284) );
  AOI22_X2 U10004 ( .A1(regBoiz_regfile_29__13_), .A2(net367001), .B1(
        regBoiz_regfile_31__13_), .B2(net366969), .ZN(n7402) );
  NOR2_X2 U10005 ( .A1(n12043), .A2(n12046), .ZN(n12044) );
  OAI21_X1 U10006 ( .B1(n5698), .B2(n7679), .A(n5093), .ZN(n7680) );
  OAI21_X1 U10007 ( .B1(n5699), .B2(n7685), .A(n5093), .ZN(n7687) );
  OAI21_X1 U10008 ( .B1(n7692), .B2(n7691), .A(n5093), .ZN(n7694) );
  OAI21_X1 U10009 ( .B1(n5451), .B2(n7700), .A(n5107), .ZN(n7702) );
  OAI21_X1 U10010 ( .B1(n7723), .B2(n7722), .A(n5107), .ZN(n7724) );
  OAI21_X1 U10011 ( .B1(n7707), .B2(n7706), .A(n5107), .ZN(n7708) );
  OAI21_X1 U10012 ( .B1(n5697), .B2(n7729), .A(n5093), .ZN(n7730) );
  OAI21_X1 U10013 ( .B1(n5452), .B2(n7713), .A(n5093), .ZN(n7715) );
  NAND2_X1 U10014 ( .A1(n6587), .A2(net376077), .ZN(n13379) );
  NAND2_X1 U10015 ( .A1(regBoiz_regfile_8__23_), .A2(net376331), .ZN(n7785) );
  NAND2_X4 U10016 ( .A1(n11248), .A2(n11247), .ZN(n11476) );
  NAND4_X2 U10017 ( .A1(n12097), .A2(n12123), .A3(n11960), .A4(n12110), .ZN(
        n12098) );
  NAND3_X4 U10018 ( .A1(n10788), .A2(n10787), .A3(n10786), .ZN(n10821) );
  OAI211_X2 U10019 ( .C1(n10785), .C2(n10816), .A(n10784), .B(n10849), .ZN(
        n10788) );
  NAND2_X1 U10020 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  NAND2_X4 U10021 ( .A1(net361802), .A2(n10917), .ZN(n10561) );
  NOR3_X2 U10022 ( .A1(n11184), .A2(n6379), .A3(n11183), .ZN(n11235) );
  NAND2_X1 U10023 ( .A1(regBoiz_regfile_4__31_), .A2(net375929), .ZN(n6286) );
  NAND2_X2 U10024 ( .A1(n6286), .A2(n6287), .ZN(n8173) );
  INV_X8 U10025 ( .A(n11989), .ZN(n11996) );
  INV_X4 U10026 ( .A(n11823), .ZN(n12043) );
  INV_X4 U10027 ( .A(n6790), .ZN(n6789) );
  INV_X2 U10028 ( .A(n6389), .ZN(n8026) );
  MUX2_X2 U10029 ( .A(regBoiz_regfile_2__16_), .B(regBoiz_regfile_10__16_), 
        .S(net369200), .Z(n7502) );
  NAND2_X4 U10030 ( .A1(n11248), .A2(n11247), .ZN(n9841) );
  NAND2_X4 U10031 ( .A1(n11647), .A2(n11646), .ZN(n11591) );
  NAND2_X4 U10032 ( .A1(n11658), .A2(n11657), .ZN(n11703) );
  NAND2_X4 U10033 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  NAND3_X4 U10034 ( .A1(n12452), .A2(n6392), .A3(n12557), .ZN(n12453) );
  NAND3_X2 U10035 ( .A1(n6993), .A2(n6793), .A3(n8144), .ZN(net364803) );
  INV_X2 U10036 ( .A(n8144), .ZN(n8138) );
  NAND3_X2 U10037 ( .A1(n8144), .A2(n8143), .A3(n8142), .ZN(n8149) );
  NOR2_X2 U10038 ( .A1(net366949), .A2(n8053), .ZN(n8049) );
  AOI21_X2 U10039 ( .B1(n10810), .B2(n10887), .A(n10809), .ZN(n10813) );
  NAND2_X4 U10040 ( .A1(n12102), .A2(n5934), .ZN(n12150) );
  NAND3_X2 U10041 ( .A1(n12151), .A2(n12150), .A3(aluBoi_multBoi_temppp[57]), 
        .ZN(n12132) );
  AOI21_X2 U10042 ( .B1(n8098), .B2(n8097), .A(net366925), .ZN(n8099) );
  AOI21_X2 U10043 ( .B1(n10550), .B2(n6003), .A(net368195), .ZN(n10555) );
  NAND2_X1 U10044 ( .A1(regBoiz_regfile_30__29_), .A2(n340), .ZN(n351) );
  INV_X8 U10045 ( .A(n11700), .ZN(n11512) );
  NAND2_X4 U10046 ( .A1(net365336), .A2(n5140), .ZN(net364941) );
  NAND2_X4 U10047 ( .A1(n11917), .A2(n11953), .ZN(n12123) );
  NAND2_X4 U10048 ( .A1(n11490), .A2(n6064), .ZN(n11421) );
  INV_X4 U10049 ( .A(n10451), .ZN(n8055) );
  NAND2_X4 U10050 ( .A1(n10567), .A2(n10568), .ZN(n10682) );
  NAND2_X4 U10051 ( .A1(n7531), .A2(net361491), .ZN(n11182) );
  OAI21_X2 U10052 ( .B1(n5675), .B2(n6736), .A(n541), .ZN(n3788) );
  OAI21_X2 U10053 ( .B1(n11831), .B2(n11830), .A(n4979), .ZN(n12011) );
  NAND2_X4 U10054 ( .A1(n8072), .A2(net366939), .ZN(n10436) );
  INV_X8 U10055 ( .A(net364904), .ZN(net364968) );
  INV_X16 U10056 ( .A(n6792), .ZN(n6782) );
  NAND2_X4 U10057 ( .A1(n11498), .A2(n11497), .ZN(n11843) );
  NAND2_X4 U10058 ( .A1(n11866), .A2(n11865), .ZN(n11864) );
  NAND2_X4 U10059 ( .A1(n11064), .A2(n11065), .ZN(n11175) );
  NAND3_X2 U10060 ( .A1(n11861), .A2(n11499), .A3(n11699), .ZN(n11504) );
  NAND2_X4 U10061 ( .A1(n6240), .A2(n12425), .ZN(n12456) );
  NAND2_X2 U10062 ( .A1(n8176), .A2(net368862), .ZN(n6288) );
  NAND2_X2 U10063 ( .A1(n8175), .A2(net366987), .ZN(n6289) );
  MUX2_X2 U10064 ( .A(n6291), .B(n6292), .S(net375727), .Z(n6290) );
  NAND2_X4 U10065 ( .A1(n12168), .A2(n12069), .ZN(n11989) );
  INV_X8 U10066 ( .A(n11300), .ZN(n11248) );
  NAND2_X4 U10067 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  INV_X16 U10068 ( .A(net368225), .ZN(net368221) );
  INV_X2 U10069 ( .A(net368225), .ZN(net368223) );
  INV_X4 U10070 ( .A(n11853), .ZN(n11866) );
  NOR2_X2 U10071 ( .A1(n11626), .A2(n11627), .ZN(n11634) );
  NAND2_X1 U10072 ( .A1(regBoiz_regfile_10__31_), .A2(net367593), .ZN(n1084)
         );
  MUX2_X1 U10073 ( .A(regBoiz_regfile_10__31_), .B(regBoiz_regfile_11__31_), 
        .S(net369157), .Z(n8331) );
  INV_X32 U10074 ( .A(net368548), .ZN(net362297) );
  INV_X8 U10075 ( .A(n5892), .ZN(n6544) );
  NAND2_X1 U10076 ( .A1(regBoiz_regfile_6__31_), .A2(net375867), .ZN(n6293) );
  NAND2_X1 U10077 ( .A1(regBoiz_regfile_14__31_), .A2(net375510), .ZN(n6294)
         );
  NAND2_X2 U10078 ( .A1(n6293), .A2(n6294), .ZN(n8172) );
  XNOR2_X1 U10079 ( .A(n10492), .B(n10491), .ZN(n10493) );
  NAND2_X4 U10080 ( .A1(n10471), .A2(n10492), .ZN(net362318) );
  XNOR2_X1 U10081 ( .A(net362224), .B(net362256), .ZN(n6441) );
  NAND2_X4 U10082 ( .A1(n10847), .A2(n10953), .ZN(n10848) );
  NAND4_X4 U10083 ( .A1(n6279), .A2(n10722), .A3(n10906), .A4(n10684), .ZN(
        n10612) );
  NOR2_X1 U10084 ( .A1(net366925), .A2(n5637), .ZN(n7678) );
  AOI21_X1 U10085 ( .B1(n7792), .B2(n7791), .A(net366925), .ZN(n7793) );
  AOI21_X1 U10086 ( .B1(n8092), .B2(n8091), .A(net366925), .ZN(n8093) );
  NOR2_X1 U10087 ( .A1(net366925), .A2(n5638), .ZN(n7462) );
  NOR2_X1 U10088 ( .A1(net366925), .A2(n5420), .ZN(n7469) );
  NOR2_X1 U10089 ( .A1(net366925), .A2(n5584), .ZN(n7470) );
  AOI21_X2 U10090 ( .B1(n8110), .B2(n8109), .A(net366925), .ZN(n8111) );
  INV_X8 U10091 ( .A(n6536), .ZN(n6537) );
  INV_X8 U10092 ( .A(n6537), .ZN(n10995) );
  OAI21_X2 U10093 ( .B1(n11513), .B2(n11512), .A(n11738), .ZN(n11514) );
  INV_X8 U10094 ( .A(n10738), .ZN(n10641) );
  NOR2_X2 U10095 ( .A1(net369316), .A2(n8122), .ZN(n8043) );
  NOR3_X2 U10096 ( .A1(n8122), .A2(n8121), .A3(net366997), .ZN(n8125) );
  XNOR2_X2 U10097 ( .A(n11779), .B(n6215), .ZN(n11755) );
  NAND2_X4 U10098 ( .A1(n11754), .A2(n11805), .ZN(n11779) );
  NAND3_X2 U10099 ( .A1(net368571), .A2(n11524), .A3(n11523), .ZN(n11605) );
  NAND2_X2 U10100 ( .A1(n11128), .A2(net369286), .ZN(n11132) );
  NAND2_X4 U10101 ( .A1(n12242), .A2(n12085), .ZN(n12243) );
  NAND2_X4 U10102 ( .A1(n6032), .A2(n12104), .ZN(n12009) );
  INV_X16 U10103 ( .A(net378321), .ZN(net366949) );
  NAND2_X4 U10104 ( .A1(net360821), .A2(n6541), .ZN(n10684) );
  NAND2_X4 U10105 ( .A1(n10684), .A2(net368211), .ZN(n10689) );
  NAND2_X4 U10106 ( .A1(n10842), .A2(n10829), .ZN(n10738) );
  NOR3_X4 U10107 ( .A1(n11859), .A2(n11858), .A3(n6092), .ZN(n11860) );
  NAND2_X2 U10108 ( .A1(n11400), .A2(n11601), .ZN(n11393) );
  INV_X8 U10109 ( .A(net366945), .ZN(net366923) );
  AOI21_X2 U10110 ( .B1(n7820), .B2(n7819), .A(net366927), .ZN(n7821) );
  NAND2_X4 U10111 ( .A1(n10837), .A2(n5870), .ZN(net362194) );
  NAND2_X2 U10112 ( .A1(n12538), .A2(net359462), .ZN(net359497) );
  OAI211_X1 U10113 ( .C1(iaddr[7]), .C2(n5385), .A(n12859), .B(n6603), .ZN(
        n12861) );
  OAI211_X1 U10114 ( .C1(iaddr[7]), .C2(n10318), .A(n12854), .B(n6603), .ZN(
        n12856) );
  OAI211_X1 U10115 ( .C1(iaddr[11]), .C2(n10264), .A(n12811), .B(n6603), .ZN(
        n12813) );
  OAI211_X1 U10116 ( .C1(iaddr[16]), .C2(n10199), .A(n12765), .B(n6603), .ZN(
        n12767) );
  OAI211_X1 U10117 ( .C1(iaddr[17]), .C2(n10186), .A(n12750), .B(n6603), .ZN(
        n12752) );
  OAI211_X1 U10118 ( .C1(iaddr[23]), .C2(n9986), .A(n12687), .B(n6603), .ZN(
        n12689) );
  OAI211_X1 U10119 ( .C1(iaddr[22]), .C2(n10122), .A(n12705), .B(n6603), .ZN(
        n12707) );
  OAI211_X1 U10120 ( .C1(iaddr[27]), .C2(n5886), .A(n12645), .B(n6603), .ZN(
        n12647) );
  INV_X2 U10121 ( .A(n12687), .ZN(n12682) );
  NAND2_X1 U10122 ( .A1(iaddr[7]), .A2(n5385), .ZN(n12859) );
  AOI21_X1 U10123 ( .B1(n10286), .B2(n12765), .A(n6434), .ZN(n10187) );
  NOR2_X1 U10124 ( .A1(n12705), .A2(n6551), .ZN(n10116) );
  NOR2_X1 U10125 ( .A1(n12645), .A2(n6551), .ZN(n10051) );
  NOR2_X1 U10126 ( .A1(n12687), .A2(n6551), .ZN(n10104) );
  AOI21_X1 U10127 ( .B1(n10286), .B2(n12750), .A(MoLanBoJ), .ZN(n10182) );
  AOI21_X1 U10128 ( .B1(n10286), .B2(n12811), .A(MoLanBoJ), .ZN(n10260) );
  NAND2_X1 U10129 ( .A1(n6571), .A2(n12705), .ZN(n10114) );
  NAND2_X1 U10130 ( .A1(n6571), .A2(n12645), .ZN(n10049) );
  NAND2_X1 U10131 ( .A1(n10318), .A2(iaddr[7]), .ZN(n12854) );
  NAND4_X4 U10132 ( .A1(iaddr[6]), .A2(iaddr[5]), .A3(iaddr[8]), .A4(iaddr[7]), 
        .ZN(n12830) );
  NAND2_X4 U10133 ( .A1(n10990), .A2(n10989), .ZN(n11046) );
  NAND2_X4 U10134 ( .A1(net362361), .A2(n10513), .ZN(n10536) );
  NOR2_X2 U10135 ( .A1(n5997), .A2(n11711), .ZN(n11652) );
  INV_X8 U10136 ( .A(n6147), .ZN(n10528) );
  OAI22_X4 U10137 ( .A1(n8032), .A2(n9850), .B1(n8031), .B2(n8030), .ZN(n10477) );
  NOR3_X2 U10138 ( .A1(n10918), .A2(n5259), .A3(net377531), .ZN(n10919) );
  INV_X2 U10139 ( .A(n12137), .ZN(n12092) );
  INV_X1 U10140 ( .A(n12418), .ZN(n12421) );
  NAND2_X4 U10141 ( .A1(n10568), .A2(n10567), .ZN(n10780) );
  NAND3_X4 U10142 ( .A1(n10835), .A2(n6435), .A3(n10856), .ZN(n10953) );
  NAND2_X4 U10143 ( .A1(net361749), .A2(net361546), .ZN(n11130) );
  INV_X2 U10144 ( .A(n10725), .ZN(n10569) );
  OAI21_X1 U10145 ( .B1(n6562), .B2(n9566), .A(net377607), .ZN(n9567) );
  OAI21_X1 U10146 ( .B1(net377607), .B2(n6564), .A(n6561), .ZN(n9564) );
  INV_X1 U10147 ( .A(n6240), .ZN(n12409) );
  NAND2_X1 U10148 ( .A1(n9377), .A2(net377607), .ZN(n9378) );
  INV_X2 U10149 ( .A(net377607), .ZN(net360360) );
  INV_X2 U10150 ( .A(net377607), .ZN(net360539) );
  INV_X2 U10151 ( .A(net377607), .ZN(net360713) );
  NOR2_X4 U10152 ( .A1(net375793), .A2(n11339), .ZN(n11340) );
  OAI22_X4 U10153 ( .A1(n10850), .A2(net368436), .B1(n11111), .B2(net368179), 
        .ZN(net361057) );
  NAND2_X4 U10154 ( .A1(n9808), .A2(n11771), .ZN(n6334) );
  INV_X1 U10155 ( .A(n6509), .ZN(n12185) );
  INV_X2 U10156 ( .A(n6509), .ZN(n12059) );
  NAND2_X1 U10157 ( .A1(net359752), .A2(n6509), .ZN(n12269) );
  MUX2_X1 U10158 ( .A(n7018), .B(n7017), .S(net366977), .Z(n7019) );
  MUX2_X2 U10159 ( .A(n6296), .B(n6297), .S(net367035), .Z(n6295) );
  INV_X8 U10160 ( .A(net367035), .ZN(net367027) );
  INV_X2 U10161 ( .A(n6298), .ZN(n6299) );
  NAND2_X1 U10162 ( .A1(regBoiz_regfile_15__6_), .A2(n6697), .ZN(n912) );
  MUX2_X2 U10163 ( .A(n7026), .B(n7025), .S(net366933), .Z(n7027) );
  INV_X2 U10164 ( .A(net375768), .ZN(net375769) );
  MUX2_X2 U10165 ( .A(n6503), .B(n6486), .S(net375527), .Z(n6301) );
  NAND2_X1 U10166 ( .A1(regBoiz_regfile_29__1_), .A2(n6751), .ZN(n427) );
  NAND2_X1 U10167 ( .A1(regBoiz_regfile_23__1_), .A2(n6730), .ZN(n629) );
  MUX2_X2 U10168 ( .A(n6341), .B(n6303), .S(net376642), .Z(n6302) );
  INV_X2 U10169 ( .A(n6304), .ZN(n6305) );
  INV_X4 U10170 ( .A(n11718), .ZN(n6375) );
  AOI21_X2 U10171 ( .B1(n11298), .B2(n11718), .A(net368211), .ZN(n11189) );
  INV_X2 U10172 ( .A(n6306), .ZN(n6307) );
  MUX2_X2 U10173 ( .A(regBoiz_regfile_20__5_), .B(regBoiz_regfile_28__5_), .S(
        net366899), .Z(n7131) );
  INV_X4 U10174 ( .A(net367035), .ZN(net375718) );
  INV_X2 U10175 ( .A(n6308), .ZN(n6309) );
  AOI21_X1 U10176 ( .B1(n7848), .B2(net366949), .A(n5159), .ZN(n7860) );
  MUX2_X1 U10177 ( .A(regBoiz_regfile_10__11_), .B(regBoiz_regfile_11__11_), 
        .S(net376222), .Z(n7330) );
  MUX2_X1 U10178 ( .A(regBoiz_regfile_26__11_), .B(regBoiz_regfile_27__11_), 
        .S(net367023), .Z(n7309) );
  NAND2_X1 U10179 ( .A1(regBoiz_regfile_27__1_), .A2(n6745), .ZN(n494) );
  MUX2_X2 U10180 ( .A(n7116), .B(n7115), .S(net366933), .Z(n7117) );
  NAND2_X2 U10181 ( .A1(n11771), .A2(n11769), .ZN(n13532) );
  MUX2_X1 U10182 ( .A(n6299), .B(n6333), .S(net368800), .Z(n7023) );
  NAND2_X1 U10183 ( .A1(regBoiz_regfile_31__6_), .A2(n6755), .ZN(n310) );
  INV_X2 U10184 ( .A(net367043), .ZN(net375738) );
  INV_X2 U10185 ( .A(n6310), .ZN(n6311) );
  INV_X2 U10186 ( .A(n6312), .ZN(n6313) );
  INV_X16 U10187 ( .A(net375618), .ZN(net369316) );
  NAND2_X1 U10188 ( .A1(regBoiz_regfile_3__4_), .A2(n6758), .ZN(n278) );
  MUX2_X2 U10189 ( .A(n7013), .B(n7014), .S(net376417), .Z(n7030) );
  MUX2_X1 U10190 ( .A(n7133), .B(n7132), .S(net378321), .Z(n7134) );
  INV_X16 U10191 ( .A(net329432), .ZN(net368571) );
  MUX2_X2 U10192 ( .A(n7028), .B(n7027), .S(net375727), .Z(n7029) );
  MUX2_X2 U10193 ( .A(n7024), .B(n7023), .S(net366977), .Z(n7025) );
  NAND2_X1 U10194 ( .A1(regBoiz_regfile_17__4_), .A2(n6704), .ZN(n847) );
  INV_X16 U10195 ( .A(net367041), .ZN(net375713) );
  MUX2_X2 U10196 ( .A(n7142), .B(n7143), .S(net375721), .Z(n7147) );
  NAND2_X1 U10197 ( .A1(regBoiz_regfile_31__2_), .A2(n6757), .ZN(n316) );
  MUX2_X1 U10198 ( .A(n7162), .B(n7161), .S(net366967), .Z(n7163) );
  OAI21_X1 U10199 ( .B1(n6562), .B2(n9596), .A(n6511), .ZN(n9597) );
  OAI21_X1 U10200 ( .B1(n6511), .B2(n6563), .A(n6560), .ZN(n9594) );
  OAI21_X2 U10201 ( .B1(n5688), .B2(n6765), .A(n210), .ZN(n3603) );
  INV_X4 U10202 ( .A(n6331), .ZN(n7101) );
  NAND2_X1 U10203 ( .A1(regBoiz_regfile_7__7_), .A2(n6774), .ZN(n138) );
  OAI21_X2 U10204 ( .B1(n5688), .B2(n6758), .A(n278), .ZN(n3601) );
  INV_X2 U10205 ( .A(n6314), .ZN(n6315) );
  NAND2_X2 U10206 ( .A1(n7091), .A2(n6786), .ZN(n6418) );
  NAND2_X1 U10207 ( .A1(regBoiz_regfile_15__8_), .A2(n6698), .ZN(n910) );
  OAI21_X2 U10208 ( .B1(n6668), .B2(n6704), .A(n847), .ZN(n3615) );
  INV_X2 U10209 ( .A(n6317), .ZN(n6318) );
  INV_X2 U10210 ( .A(n6319), .ZN(n6320) );
  INV_X2 U10211 ( .A(n6321), .ZN(n6322) );
  NAND2_X1 U10212 ( .A1(regBoiz_regfile_13__7_), .A2(n6690), .ZN(n978) );
  INV_X2 U10213 ( .A(n6323), .ZN(n6324) );
  NAND2_X1 U10214 ( .A1(n6693), .A2(regBoiz_regfile_14__7_), .ZN(n945) );
  NAND2_X1 U10215 ( .A1(regBoiz_regfile_6__4_), .A2(n6769), .ZN(n176) );
  MUX2_X2 U10216 ( .A(n6305), .B(n6339), .S(n4978), .Z(n7096) );
  MUX2_X2 U10217 ( .A(regBoiz_regfile_6__4_), .B(regBoiz_regfile_7__4_), .S(
        net369147), .Z(n9311) );
  MUX2_X2 U10218 ( .A(n6443), .B(n6326), .S(net375867), .Z(n6325) );
  NAND2_X2 U10219 ( .A1(n7307), .A2(n6221), .ZN(n6327) );
  INV_X2 U10220 ( .A(n6329), .ZN(n6330) );
  NAND2_X1 U10221 ( .A1(regBoiz_regfile_28__10_), .A2(n6748), .ZN(n470) );
  NAND2_X1 U10222 ( .A1(regBoiz_regfile_22__10_), .A2(n6727), .ZN(n673) );
  MUX2_X2 U10223 ( .A(n6469), .B(n6340), .S(net376642), .Z(n6331) );
  MUX2_X1 U10224 ( .A(n7102), .B(n7101), .S(net366979), .Z(n7103) );
  INV_X2 U10225 ( .A(n6332), .ZN(n6333) );
  AOI21_X1 U10226 ( .B1(n9877), .B2(n6793), .A(net367019), .ZN(n9879) );
  MUX2_X1 U10227 ( .A(regBoiz_regfile_18__11_), .B(regBoiz_regfile_19__11_), 
        .S(net376223), .Z(n7327) );
  NAND2_X4 U10228 ( .A1(n11727), .A2(n6335), .ZN(n9809) );
  NAND2_X1 U10229 ( .A1(regBoiz_regfile_31__1_), .A2(n6757), .ZN(n327) );
  NOR2_X2 U10230 ( .A1(n9807), .A2(n9806), .ZN(n9808) );
  NAND2_X1 U10231 ( .A1(net376331), .A2(net367005), .ZN(n8150) );
  MUX2_X2 U10232 ( .A(regBoiz_regfile_1__9_), .B(n6407), .S(net366899), .Z(
        n7254) );
  MUX2_X1 U10233 ( .A(regBoiz_regfile_2__4_), .B(n6318), .S(net376077), .Z(
        n7094) );
  INV_X2 U10234 ( .A(n6336), .ZN(n6337) );
  INV_X2 U10235 ( .A(n6338), .ZN(n6339) );
  MUX2_X2 U10236 ( .A(n7273), .B(n7274), .S(net375618), .Z(n7275) );
  NAND2_X1 U10237 ( .A1(regBoiz_regfile_21__9_), .A2(n6724), .ZN(n676) );
  NAND2_X2 U10238 ( .A1(n7260), .A2(net375614), .ZN(n6342) );
  NAND2_X1 U10239 ( .A1(n7259), .A2(net375738), .ZN(n6343) );
  NAND2_X2 U10240 ( .A1(n6342), .A2(n6343), .ZN(n7276) );
  NAND2_X2 U10241 ( .A1(n7266), .A2(net376387), .ZN(n6344) );
  NAND2_X1 U10242 ( .A1(n7265), .A2(net378321), .ZN(n6345) );
  NAND2_X2 U10243 ( .A1(n6344), .A2(n6345), .ZN(n7274) );
  MUX2_X2 U10244 ( .A(n6347), .B(n6348), .S(net377464), .Z(n6346) );
  MUX2_X2 U10245 ( .A(n7272), .B(n7271), .S(net378321), .Z(n7273) );
  NAND2_X2 U10246 ( .A1(n7108), .A2(net375547), .ZN(n6349) );
  NAND2_X1 U10247 ( .A1(n7107), .A2(net366967), .ZN(n6350) );
  NAND2_X2 U10248 ( .A1(n6349), .A2(n6350), .ZN(n7112) );
  MUX2_X2 U10249 ( .A(n6352), .B(n6353), .S(n5245), .Z(n6351) );
  INV_X32 U10250 ( .A(net375309), .ZN(net375310) );
  NAND3_X2 U10251 ( .A1(n11113), .A2(n11105), .A3(n11106), .ZN(n11108) );
  NAND2_X1 U10252 ( .A1(regBoiz_regfile_6__26_), .A2(net376541), .ZN(n6354) );
  NAND2_X1 U10253 ( .A1(regBoiz_regfile_14__26_), .A2(net376063), .ZN(n6355)
         );
  NAND2_X2 U10254 ( .A1(n6354), .A2(n6355), .ZN(n7963) );
  NAND2_X2 U10255 ( .A1(n7964), .A2(net375547), .ZN(n6356) );
  NAND2_X1 U10256 ( .A1(n7963), .A2(net366973), .ZN(n6357) );
  NAND2_X2 U10257 ( .A1(n6356), .A2(n6357), .ZN(n7965) );
  NAND2_X2 U10258 ( .A1(n11506), .A2(n11505), .ZN(n11563) );
  OR2_X4 U10259 ( .A1(n12046), .A2(n5911), .ZN(n12049) );
  NAND2_X4 U10260 ( .A1(n11995), .A2(n5966), .ZN(n12167) );
  NOR2_X4 U10261 ( .A1(n9883), .A2(n9882), .ZN(n6358) );
  NOR2_X4 U10262 ( .A1(n9884), .A2(n6359), .ZN(n9885) );
  INV_X4 U10263 ( .A(n6358), .ZN(n6359) );
  NAND2_X2 U10264 ( .A1(n7775), .A2(n6230), .ZN(n6360) );
  NAND2_X1 U10265 ( .A1(n7774), .A2(n6788), .ZN(n6361) );
  NAND2_X2 U10266 ( .A1(n6360), .A2(n6361), .ZN(n9884) );
  NAND2_X2 U10267 ( .A1(n9884), .A2(net375929), .ZN(n6415) );
  INV_X16 U10268 ( .A(net369208), .ZN(net369202) );
  INV_X2 U10269 ( .A(n6371), .ZN(n7989) );
  INV_X8 U10270 ( .A(net368903), .ZN(net369208) );
  NAND3_X2 U10271 ( .A1(n6067), .A2(n11230), .A3(n10896), .ZN(n10901) );
  NAND2_X4 U10272 ( .A1(n12042), .A2(n12167), .ZN(n12173) );
  MUX2_X2 U10273 ( .A(regBoiz_regfile_26__26_), .B(regBoiz_regfile_18__26_), 
        .S(net369206), .Z(n7931) );
  NAND2_X4 U10274 ( .A1(n12173), .A2(n12172), .ZN(n12046) );
  NAND2_X4 U10275 ( .A1(n11668), .A2(aluBoi_multBoi_temppp[48]), .ZN(net359916) );
  MUX2_X2 U10276 ( .A(n6363), .B(n6364), .S(net369206), .Z(n6362) );
  NAND2_X2 U10277 ( .A1(n7800), .A2(net375547), .ZN(n6365) );
  NAND2_X1 U10278 ( .A1(n7799), .A2(net366973), .ZN(n6366) );
  NAND2_X2 U10279 ( .A1(n6365), .A2(n6366), .ZN(n7801) );
  MUX2_X2 U10280 ( .A(n6368), .B(n6369), .S(net366885), .Z(n6367) );
  NAND2_X1 U10281 ( .A1(regBoiz_regfile_23__23_), .A2(n6730), .ZN(n625) );
  MUX2_X1 U10282 ( .A(regBoiz_regfile_19__23_), .B(regBoiz_regfile_23__23_), 
        .S(net378321), .Z(n7772) );
  NAND3_X2 U10283 ( .A1(n10718), .A2(n10717), .A3(n10716), .ZN(n10736) );
  NAND2_X4 U10284 ( .A1(n10694), .A2(n10693), .ZN(n10845) );
  NAND3_X2 U10285 ( .A1(n7651), .A2(n7650), .A3(n7649), .ZN(n7677) );
  NOR2_X4 U10286 ( .A1(n6420), .A2(n6375), .ZN(n6374) );
  INV_X4 U10287 ( .A(n6374), .ZN(n11767) );
  NAND2_X4 U10288 ( .A1(n11520), .A2(n11519), .ZN(n6420) );
  NAND2_X4 U10289 ( .A1(n10952), .A2(net361629), .ZN(n10836) );
  NAND2_X1 U10290 ( .A1(regBoiz_regfile_12__23_), .A2(net368781), .ZN(n7783)
         );
  MUX2_X2 U10291 ( .A(n7988), .B(n7989), .S(net366999), .Z(n7993) );
  INV_X8 U10292 ( .A(net367007), .ZN(net366999) );
  OAI21_X2 U10293 ( .B1(n5683), .B2(net367593), .A(n1084), .ZN(n4499) );
  NAND2_X4 U10294 ( .A1(n11403), .A2(n6026), .ZN(n11468) );
  NAND3_X2 U10295 ( .A1(n11198), .A2(n11197), .A3(n11196), .ZN(n11201) );
  INV_X8 U10296 ( .A(n11004), .ZN(n11196) );
  NAND2_X4 U10297 ( .A1(n12262), .A2(n12261), .ZN(n12260) );
  INV_X4 U10298 ( .A(n6381), .ZN(n7799) );
  OAI22_X1 U10299 ( .A1(n7383), .A2(net367031), .B1(n7382), .B2(net367041), 
        .ZN(n7384) );
  AOI22_X2 U10300 ( .A1(regBoiz_regfile_4__13_), .A2(net367003), .B1(
        regBoiz_regfile_6__13_), .B2(net366985), .ZN(n7383) );
  INV_X2 U10301 ( .A(n6377), .ZN(n6378) );
  INV_X4 U10302 ( .A(net367027), .ZN(net375506) );
  NAND2_X2 U10303 ( .A1(n12381), .A2(n12422), .ZN(n12400) );
  NAND2_X4 U10304 ( .A1(n11151), .A2(n11150), .ZN(n11163) );
  NAND4_X4 U10305 ( .A1(n11305), .A2(n11304), .A3(n11307), .A4(n11306), .ZN(
        n11483) );
  NAND2_X4 U10306 ( .A1(n5948), .A2(n11478), .ZN(n11723) );
  NAND2_X4 U10307 ( .A1(n9828), .A2(n11191), .ZN(n11300) );
  INV_X1 U10308 ( .A(n6536), .ZN(n6379) );
  NAND2_X4 U10309 ( .A1(net361903), .A2(net378405), .ZN(net361902) );
  NAND3_X1 U10310 ( .A1(n12262), .A2(n12261), .A3(n12568), .ZN(n12267) );
  NOR2_X2 U10311 ( .A1(n5971), .A2(n12348), .ZN(n12352) );
  NOR2_X4 U10312 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  MUX2_X1 U10313 ( .A(n7453), .B(n7452), .S(net378488), .Z(n7454) );
  INV_X2 U10314 ( .A(n10536), .ZN(n10467) );
  AOI21_X1 U10315 ( .B1(n12209), .B2(net345751), .A(aluBoi_multBoi_temppp[29]), 
        .ZN(n12210) );
  NOR2_X1 U10316 ( .A1(net345751), .A2(net368209), .ZN(n10522) );
  NOR2_X2 U10317 ( .A1(net345751), .A2(net368498), .ZN(n10474) );
  AOI21_X1 U10318 ( .B1(n9684), .B2(net345751), .A(n9683), .ZN(n9685) );
  OAI21_X1 U10319 ( .B1(n6019), .B2(n9677), .A(net345751), .ZN(n8713) );
  NOR2_X2 U10320 ( .A1(n12210), .A2(n10494), .ZN(n12212) );
  OAI21_X2 U10321 ( .B1(n6565), .B2(n9678), .A(n8713), .ZN(n9085) );
  NAND2_X4 U10322 ( .A1(aluBoi_multBoi_temppp[54]), .A2(net360253), .ZN(
        net360011) );
  NOR3_X2 U10323 ( .A1(n10629), .A2(net362047), .A3(net362048), .ZN(n10630) );
  NAND2_X4 U10324 ( .A1(n10779), .A2(n10778), .ZN(n10893) );
  NAND2_X4 U10325 ( .A1(n10893), .A2(n11181), .ZN(n10913) );
  MUX2_X2 U10326 ( .A(n6382), .B(n6383), .S(net366901), .Z(n6381) );
  NOR2_X2 U10327 ( .A1(n6092), .A2(n11660), .ZN(n11499) );
  NOR2_X2 U10328 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  NAND4_X2 U10329 ( .A1(n11245), .A2(n5241), .A3(n11243), .A4(n11242), .ZN(
        n11246) );
  NAND2_X4 U10330 ( .A1(n11577), .A2(n11657), .ZN(n11850) );
  INV_X2 U10331 ( .A(n8031), .ZN(n7983) );
  NAND2_X4 U10332 ( .A1(net362256), .A2(net362224), .ZN(n10501) );
  INV_X1 U10333 ( .A(n10995), .ZN(n6384) );
  INV_X2 U10334 ( .A(net361278), .ZN(net361326) );
  AOI21_X2 U10335 ( .B1(n7618), .B2(n7617), .A(net366967), .ZN(n7621) );
  AOI21_X2 U10336 ( .B1(regBoiz_regfile_16__19_), .B2(net366949), .A(n6793), 
        .ZN(n7618) );
  NAND2_X1 U10337 ( .A1(regBoiz_regfile_20__19_), .A2(net366919), .ZN(n7617)
         );
  OAI211_X1 U10338 ( .C1(net366933), .C2(n5582), .A(n6794), .B(n7619), .ZN(
        n7620) );
  NOR3_X2 U10339 ( .A1(n11000), .A2(net375435), .A3(n6194), .ZN(n10774) );
  OAI21_X4 U10340 ( .B1(n12098), .B2(n12099), .A(n6033), .ZN(n12135) );
  AOI21_X4 U10341 ( .B1(n11272), .B2(n11460), .A(n11270), .ZN(n11273) );
  NAND3_X2 U10342 ( .A1(n11816), .A2(n11820), .A3(n11815), .ZN(n6385) );
  NAND2_X4 U10343 ( .A1(n11806), .A2(n11807), .ZN(n11816) );
  AOI21_X2 U10344 ( .B1(regBoiz_regfile_2__19_), .B2(net366949), .A(n6782), 
        .ZN(n7615) );
  AOI21_X2 U10345 ( .B1(n7824), .B2(n7823), .A(net366949), .ZN(n7828) );
  NAND2_X4 U10346 ( .A1(n11750), .A2(n11584), .ZN(n11870) );
  INV_X2 U10347 ( .A(n10619), .ZN(n6387) );
  INV_X8 U10348 ( .A(n13526), .ZN(n6514) );
  INV_X16 U10349 ( .A(n6515), .ZN(n12053) );
  INV_X8 U10350 ( .A(n9897), .ZN(n11245) );
  NAND2_X1 U10351 ( .A1(net359766), .A2(net359767), .ZN(n12337) );
  NAND2_X1 U10352 ( .A1(n11213), .A2(n11214), .ZN(n11283) );
  NAND2_X4 U10353 ( .A1(n11214), .A2(n11213), .ZN(n11376) );
  OAI22_X2 U10354 ( .A1(n12060), .A2(net368462), .B1(n6049), .B2(net368195), 
        .ZN(n12176) );
  NOR2_X4 U10355 ( .A1(n11319), .A2(net361090), .ZN(n11320) );
  INV_X8 U10356 ( .A(net361053), .ZN(net361090) );
  NAND2_X4 U10357 ( .A1(n11503), .A2(n11502), .ZN(n11577) );
  OAI211_X4 U10358 ( .C1(n8059), .C2(n8058), .A(n8056), .B(n8057), .ZN(n8060)
         );
  INV_X32 U10359 ( .A(net376602), .ZN(net361801) );
  NAND2_X4 U10360 ( .A1(n10454), .A2(n6075), .ZN(net334218) );
  AOI22_X4 U10361 ( .A1(n10472), .A2(n6388), .B1(net375435), .B2(n10472), .ZN(
        net375434) );
  AND2_X2 U10362 ( .A1(n6251), .A2(n10473), .ZN(n6388) );
  OAI211_X1 U10363 ( .C1(net360583), .C2(n11697), .A(n12225), .B(net100619), 
        .ZN(n11698) );
  NAND2_X4 U10364 ( .A1(n6787), .A2(net375650), .ZN(n7943) );
  INV_X1 U10365 ( .A(n7943), .ZN(n7935) );
  NOR3_X2 U10366 ( .A1(n7943), .A2(net366919), .A3(net366997), .ZN(n7933) );
  INV_X2 U10367 ( .A(net362158), .ZN(net362157) );
  NAND2_X4 U10368 ( .A1(n11149), .A2(net361292), .ZN(n11160) );
  OAI21_X4 U10369 ( .B1(n11629), .B2(n11630), .A(n6552), .ZN(n11633) );
  NAND2_X4 U10370 ( .A1(n12456), .A2(n12557), .ZN(n12454) );
  MUX2_X2 U10371 ( .A(n6390), .B(n6391), .S(n6790), .Z(n6389) );
  OAI21_X4 U10372 ( .B1(n12395), .B2(n6123), .A(n12401), .ZN(n12396) );
  INV_X8 U10373 ( .A(n12016), .ZN(n11792) );
  NAND2_X4 U10374 ( .A1(net362230), .A2(net362229), .ZN(n10535) );
  NAND4_X1 U10375 ( .A1(n10959), .A2(n10856), .A3(n10957), .A4(n11042), .ZN(
        n10960) );
  NAND2_X4 U10376 ( .A1(net361802), .A2(net361801), .ZN(n10696) );
  NAND2_X4 U10377 ( .A1(n10609), .A2(n6543), .ZN(n10746) );
  INV_X4 U10378 ( .A(n11825), .ZN(n11818) );
  NAND3_X2 U10379 ( .A1(n11816), .A2(n11820), .A3(n11815), .ZN(n11825) );
  INV_X8 U10380 ( .A(n12451), .ZN(n12373) );
  NAND3_X4 U10381 ( .A1(n11081), .A2(n11080), .A3(n6094), .ZN(n11324) );
  OAI21_X2 U10382 ( .B1(net378128), .B2(n11034), .A(n10961), .ZN(n10962) );
  NAND2_X1 U10383 ( .A1(regBoiz_regfile_25__10_), .A2(n6738), .ZN(n571) );
  NAND2_X1 U10384 ( .A1(regBoiz_regfile_19__10_), .A2(n6712), .ZN(n805) );
  INV_X8 U10385 ( .A(net367007), .ZN(net367005) );
  INV_X8 U10386 ( .A(net367011), .ZN(net366991) );
  INV_X2 U10387 ( .A(n6395), .ZN(n6396) );
  MUX2_X1 U10388 ( .A(n7281), .B(n7280), .S(net366981), .Z(n7282) );
  MUX2_X2 U10389 ( .A(n7303), .B(n7302), .S(net366927), .Z(n7304) );
  NAND3_X2 U10390 ( .A1(n10608), .A2(n10607), .A3(n10606), .ZN(n10609) );
  OAI21_X2 U10391 ( .B1(n5649), .B2(n6747), .A(n470), .ZN(n3824) );
  NOR2_X2 U10392 ( .A1(n12041), .A2(n12040), .ZN(n12045) );
  OAI21_X2 U10393 ( .B1(n5649), .B2(n6725), .A(n673), .ZN(n3818) );
  NAND2_X1 U10394 ( .A1(regBoiz_regfile_26__10_), .A2(n6742), .ZN(n538) );
  NAND3_X2 U10395 ( .A1(n10919), .A2(n10920), .A3(n10921), .ZN(n10922) );
  INV_X16 U10396 ( .A(n13529), .ZN(n6538) );
  NAND3_X4 U10397 ( .A1(n7960), .A2(n7961), .A3(n7962), .ZN(n9788) );
  NAND2_X4 U10398 ( .A1(n10683), .A2(net361984), .ZN(n10889) );
  INV_X8 U10399 ( .A(n6428), .ZN(n12464) );
  NOR2_X1 U10400 ( .A1(n5989), .A2(n6428), .ZN(n12200) );
  NAND2_X1 U10401 ( .A1(n12464), .A2(n12359), .ZN(n12075) );
  NAND2_X2 U10402 ( .A1(n7287), .A2(net375547), .ZN(n6401) );
  NAND2_X1 U10403 ( .A1(n7286), .A2(net366979), .ZN(n6402) );
  NAND2_X2 U10404 ( .A1(n6401), .A2(n6402), .ZN(n7288) );
  MUX2_X2 U10405 ( .A(n7289), .B(n7288), .S(net366927), .Z(n7290) );
  MUX2_X2 U10406 ( .A(n6404), .B(n6405), .S(net376417), .Z(n6403) );
  INV_X2 U10407 ( .A(n6406), .ZN(n6407) );
  MUX2_X2 U10408 ( .A(n7256), .B(n7255), .S(net366981), .Z(n7257) );
  NAND2_X4 U10409 ( .A1(n12449), .A2(n6113), .ZN(n12425) );
  INV_X8 U10410 ( .A(n12394), .ZN(n12368) );
  MUX2_X2 U10411 ( .A(n7264), .B(n7263), .S(net366981), .Z(n7265) );
  NAND2_X4 U10412 ( .A1(net364968), .A2(daddr[8]), .ZN(n10703) );
  NAND2_X4 U10413 ( .A1(net366939), .A2(net367043), .ZN(n8031) );
  INV_X1 U10414 ( .A(net362256), .ZN(net375336) );
  NOR4_X4 U10415 ( .A1(net364968), .A2(n8053), .A3(net366933), .A4(n8052), 
        .ZN(n8054) );
  MUX2_X1 U10416 ( .A(n7258), .B(n7257), .S(net378321), .Z(n7259) );
  INV_X8 U10417 ( .A(n12423), .ZN(n12392) );
  OAI21_X4 U10418 ( .B1(n12366), .B2(n12429), .A(n12365), .ZN(n12367) );
  NAND2_X4 U10419 ( .A1(n10640), .A2(n10714), .ZN(n10829) );
  INV_X4 U10420 ( .A(n10840), .ZN(n10640) );
  NAND2_X4 U10421 ( .A1(n8024), .A2(n8023), .ZN(n10475) );
  OAI21_X2 U10422 ( .B1(n10435), .B2(net366921), .A(n5972), .ZN(n8059) );
  OAI21_X2 U10423 ( .B1(net368201), .B2(n10461), .A(n10573), .ZN(n10462) );
  NAND2_X4 U10424 ( .A1(n11784), .A2(net360474), .ZN(n11867) );
  INV_X8 U10425 ( .A(n11809), .ZN(n11821) );
  OAI21_X4 U10426 ( .B1(n6428), .B2(n12435), .A(n12357), .ZN(n12191) );
  INV_X2 U10427 ( .A(net361512), .ZN(net361509) );
  NAND2_X1 U10428 ( .A1(n10924), .A2(net368195), .ZN(n10925) );
  NAND2_X1 U10429 ( .A1(n10924), .A2(n6539), .ZN(n10923) );
  NAND2_X4 U10430 ( .A1(n11386), .A2(n11385), .ZN(n11641) );
  NAND2_X2 U10431 ( .A1(n9842), .A2(n9845), .ZN(n13535) );
  NAND3_X2 U10432 ( .A1(n11236), .A2(n11235), .A3(n11237), .ZN(n11186) );
  INV_X8 U10433 ( .A(n11282), .ZN(n11403) );
  INV_X8 U10434 ( .A(n6420), .ZN(n6518) );
  INV_X8 U10435 ( .A(net375279), .ZN(net375309) );
  NOR2_X1 U10436 ( .A1(net376331), .A2(n6782), .ZN(n7336) );
  NAND2_X1 U10437 ( .A1(n10644), .A2(n6282), .ZN(net362028) );
  INV_X16 U10438 ( .A(n6552), .ZN(n6553) );
  NAND2_X4 U10439 ( .A1(n11512), .A2(n11738), .ZN(n11854) );
  INV_X8 U10440 ( .A(n8106), .ZN(n7670) );
  NAND3_X2 U10441 ( .A1(n11196), .A2(n11060), .A3(n11061), .ZN(n11063) );
  AOI22_X4 U10442 ( .A1(net360821), .A2(n10579), .B1(n10485), .B2(net368498), 
        .ZN(n10540) );
  NAND4_X2 U10443 ( .A1(n10484), .A2(n10483), .A3(net362256), .A4(n10570), 
        .ZN(n10487) );
  NAND2_X4 U10444 ( .A1(net368215), .A2(n10482), .ZN(n10483) );
  NAND2_X4 U10445 ( .A1(n8178), .A2(n8179), .ZN(n8182) );
  NAND2_X1 U10446 ( .A1(n12392), .A2(n12243), .ZN(n12038) );
  XNOR2_X1 U10447 ( .A(n5274), .B(n11427), .ZN(n11314) );
  NAND3_X4 U10448 ( .A1(n11466), .A2(n11627), .A3(n11465), .ZN(n11647) );
  INV_X32 U10449 ( .A(net366935), .ZN(net366947) );
  NAND2_X4 U10450 ( .A1(n10607), .A2(net361801), .ZN(n10929) );
  NAND3_X2 U10451 ( .A1(n10438), .A2(net369316), .A3(n10439), .ZN(n10440) );
  NAND2_X4 U10452 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  NAND3_X2 U10453 ( .A1(n10723), .A2(n11232), .A3(n11242), .ZN(n11233) );
  NAND3_X2 U10454 ( .A1(n11242), .A2(n10906), .A3(n11232), .ZN(n11608) );
  NAND2_X4 U10455 ( .A1(n10552), .A2(n10551), .ZN(n10553) );
  NAND4_X2 U10456 ( .A1(n11042), .A2(n10957), .A3(n10958), .A4(n10839), .ZN(
        n10830) );
  NAND2_X4 U10457 ( .A1(n12451), .A2(n5937), .ZN(n12237) );
  NAND2_X4 U10458 ( .A1(n5896), .A2(n6063), .ZN(n11453) );
  NOR2_X1 U10459 ( .A1(n12292), .A2(n12291), .ZN(n12295) );
  INV_X8 U10460 ( .A(n11590), .ZN(n11798) );
  NAND2_X4 U10461 ( .A1(n11589), .A2(n11639), .ZN(n11590) );
  NAND3_X2 U10462 ( .A1(n10780), .A2(n5952), .A3(net361984), .ZN(n11231) );
  NAND2_X1 U10463 ( .A1(net361356), .A2(net376121), .ZN(n11142) );
  NAND2_X4 U10464 ( .A1(n11981), .A2(n6419), .ZN(n12204) );
  OAI21_X2 U10465 ( .B1(n5675), .B2(n6722), .A(n676), .ZN(n3784) );
  NOR2_X1 U10466 ( .A1(net364882), .A2(n5944), .ZN(n8126) );
  OAI21_X4 U10467 ( .B1(n10555), .B2(n10554), .A(n10553), .ZN(n10559) );
  AOI21_X1 U10468 ( .B1(n12233), .B2(n12232), .A(n12240), .ZN(n12234) );
  NAND2_X4 U10469 ( .A1(n11791), .A2(n11790), .ZN(n12016) );
  INV_X8 U10470 ( .A(n10697), .ZN(n10782) );
  NOR3_X2 U10471 ( .A1(n11950), .A2(n11949), .A3(n11948), .ZN(n11958) );
  NAND2_X4 U10472 ( .A1(n11876), .A2(n11999), .ZN(n12015) );
  INV_X16 U10473 ( .A(n6518), .ZN(n6519) );
  INV_X8 U10474 ( .A(n10929), .ZN(n11230) );
  NAND3_X2 U10475 ( .A1(n6046), .A2(n10588), .A3(n10587), .ZN(net361890) );
  XNOR2_X1 U10476 ( .A(n6097), .B(n11989), .ZN(n11985) );
  NAND2_X4 U10477 ( .A1(n11785), .A2(n11786), .ZN(n11809) );
  NAND3_X2 U10478 ( .A1(n12406), .A2(n12407), .A3(n12405), .ZN(n12413) );
  NAND3_X4 U10479 ( .A1(n12268), .A2(n12267), .A3(n12266), .ZN(n12426) );
  NOR2_X4 U10480 ( .A1(n10972), .A2(n10904), .ZN(n10911) );
  NAND3_X2 U10481 ( .A1(n11734), .A2(n11420), .A3(n11418), .ZN(n11419) );
  NAND3_X2 U10482 ( .A1(n11423), .A2(n11424), .A3(n11422), .ZN(n11439) );
  NAND2_X4 U10483 ( .A1(daddr[5]), .A2(net362342), .ZN(n10562) );
  NAND2_X4 U10484 ( .A1(net361491), .A2(n7379), .ZN(n9812) );
  NAND2_X4 U10485 ( .A1(net362231), .A2(n10534), .ZN(net362050) );
  OAI21_X2 U10486 ( .B1(n6251), .B2(net375336), .A(n10485), .ZN(n10539) );
  NAND2_X4 U10487 ( .A1(n12188), .A2(n12254), .ZN(n12278) );
  NAND2_X4 U10488 ( .A1(n11377), .A2(n11401), .ZN(n11597) );
  NAND2_X4 U10489 ( .A1(n11632), .A2(n11631), .ZN(n11824) );
  NAND4_X1 U10490 ( .A1(net368215), .A2(net362361), .A3(net362224), .A4(n5956), 
        .ZN(n10459) );
  NAND2_X2 U10491 ( .A1(n8028), .A2(net366979), .ZN(n6411) );
  NAND2_X2 U10492 ( .A1(n8029), .A2(net375547), .ZN(n6412) );
  NAND2_X2 U10493 ( .A1(n6411), .A2(n6412), .ZN(n8030) );
  INV_X4 U10494 ( .A(n6413), .ZN(n6414) );
  NAND2_X1 U10495 ( .A1(n11624), .A2(n11400), .ZN(n11277) );
  INV_X8 U10496 ( .A(n11624), .ZN(n11271) );
  NAND2_X1 U10497 ( .A1(n9881), .A2(net376374), .ZN(n6416) );
  NAND2_X2 U10498 ( .A1(n6415), .A2(n6416), .ZN(n7782) );
  NAND2_X4 U10499 ( .A1(n12368), .A2(n12384), .ZN(n12376) );
  NAND2_X4 U10500 ( .A1(n11681), .A2(aluBoi_multBoi_temppp[50]), .ZN(net360266) );
  NAND3_X2 U10501 ( .A1(n11245), .A2(n11244), .A3(n5929), .ZN(n11004) );
  NAND2_X4 U10502 ( .A1(n11845), .A2(n11868), .ZN(n11884) );
  NAND2_X4 U10503 ( .A1(n12447), .A2(n12446), .ZN(n12557) );
  XNOR2_X2 U10504 ( .A(n6419), .B(n6511), .ZN(n12248) );
  NAND2_X2 U10505 ( .A1(n11936), .A2(n11935), .ZN(n11942) );
  NAND2_X1 U10506 ( .A1(n12244), .A2(n12245), .ZN(n12159) );
  OAI22_X1 U10507 ( .A1(n10101), .A2(net368446), .B1(net368187), .B2(n11833), 
        .ZN(n11790) );
  OAI21_X1 U10508 ( .B1(n5878), .B2(net368179), .A(n12458), .ZN(n12583) );
  NAND2_X1 U10509 ( .A1(n12250), .A2(n12252), .ZN(n12354) );
  NAND2_X4 U10510 ( .A1(n12253), .A2(n12252), .ZN(n12573) );
  INV_X8 U10511 ( .A(n6796), .ZN(n6794) );
  NAND2_X4 U10512 ( .A1(net360904), .A2(net377611), .ZN(n10551) );
  NAND2_X4 U10513 ( .A1(net362270), .A2(net362297), .ZN(net362179) );
  INV_X16 U10514 ( .A(net366937), .ZN(net366951) );
  NAND2_X4 U10515 ( .A1(n10888), .A2(n11094), .ZN(net361524) );
  OAI21_X4 U10516 ( .B1(n12330), .B2(net359540), .A(net377689), .ZN(n11697) );
  XNOR2_X2 U10517 ( .A(n5029), .B(aluBoi_multBoi_temppp[41]), .ZN(net369197)
         );
  NAND3_X2 U10518 ( .A1(n11334), .A2(n11333), .A3(n11740), .ZN(n11276) );
  NAND2_X4 U10519 ( .A1(n11944), .A2(n11920), .ZN(n11946) );
  OAI21_X2 U10520 ( .B1(n10528), .B2(n5002), .A(net362297), .ZN(n8700) );
  AOI21_X2 U10521 ( .B1(n12436), .B2(n6399), .A(n12466), .ZN(n12439) );
  NAND2_X4 U10522 ( .A1(n12202), .A2(n12201), .ZN(n12233) );
  NAND3_X2 U10523 ( .A1(n12018), .A2(n5888), .A3(n12200), .ZN(n12201) );
  OAI21_X2 U10524 ( .B1(n12373), .B2(n12372), .A(n12425), .ZN(n12374) );
  NOR2_X4 U10525 ( .A1(n11570), .A2(n11569), .ZN(n11544) );
  NAND2_X4 U10526 ( .A1(net361491), .A2(n7456), .ZN(n9843) );
  NAND2_X4 U10527 ( .A1(n11308), .A2(n11309), .ZN(n11385) );
  NAND2_X4 U10528 ( .A1(n10537), .A2(net368501), .ZN(n11296) );
  NAND2_X2 U10529 ( .A1(n12465), .A2(n6139), .ZN(n12364) );
  INV_X8 U10530 ( .A(n8060), .ZN(n10454) );
  NAND2_X4 U10531 ( .A1(n5006), .A2(n11900), .ZN(n11907) );
  NAND2_X2 U10532 ( .A1(n12528), .A2(n12336), .ZN(net359756) );
  INV_X2 U10533 ( .A(n12406), .ZN(n12304) );
  NAND3_X2 U10534 ( .A1(n12005), .A2(n12004), .A3(n5943), .ZN(n12006) );
  NOR2_X2 U10535 ( .A1(n10955), .A2(n10824), .ZN(n10825) );
  NAND2_X4 U10536 ( .A1(n11452), .A2(n11687), .ZN(n11664) );
  INV_X2 U10537 ( .A(n12135), .ZN(n12102) );
  NAND2_X1 U10538 ( .A1(n11894), .A2(n11895), .ZN(n11915) );
  NAND2_X2 U10539 ( .A1(n7092), .A2(n6221), .ZN(n6417) );
  NAND2_X2 U10540 ( .A1(n6417), .A2(n6418), .ZN(n7093) );
  INV_X1 U10541 ( .A(n12182), .ZN(n6421) );
  NAND2_X4 U10542 ( .A1(n12303), .A2(net129670), .ZN(net359462) );
  NOR2_X2 U10543 ( .A1(n12508), .A2(net360265), .ZN(net360278) );
  NAND3_X2 U10544 ( .A1(n11879), .A2(n11878), .A3(n11880), .ZN(n11997) );
  INV_X1 U10545 ( .A(n6004), .ZN(n12379) );
  OAI21_X4 U10546 ( .B1(n12384), .B2(n12385), .A(n6240), .ZN(n12415) );
  XOR2_X2 U10547 ( .A(n10795), .B(n10794), .Z(n6429) );
  NAND3_X2 U10548 ( .A1(n6071), .A2(n11129), .A3(n11130), .ZN(n11100) );
  NOR3_X1 U10549 ( .A1(n12337), .A2(net359513), .A3(n6053), .ZN(n12338) );
  INV_X1 U10550 ( .A(net359481), .ZN(net359673) );
  NOR2_X2 U10551 ( .A1(n11031), .A2(n11032), .ZN(n11033) );
  AOI21_X2 U10552 ( .B1(n11945), .B2(net360235), .A(n11920), .ZN(n11926) );
  NAND2_X2 U10553 ( .A1(aluBoi_multBoi_temppp[52]), .A2(net360235), .ZN(n11938) );
  NAND2_X4 U10554 ( .A1(n6085), .A2(n11835), .ZN(net360235) );
  NAND3_X2 U10555 ( .A1(n11855), .A2(n11849), .A3(n11850), .ZN(n11758) );
  NAND2_X4 U10556 ( .A1(n11434), .A2(n11433), .ZN(net360620) );
  NAND2_X4 U10557 ( .A1(net362253), .A2(net368548), .ZN(n10526) );
  NAND3_X2 U10558 ( .A1(n12031), .A2(n12123), .A3(n11566), .ZN(n11940) );
  NAND2_X4 U10559 ( .A1(n11329), .A2(n11328), .ZN(n11547) );
  NAND2_X4 U10560 ( .A1(net361073), .A2(n11327), .ZN(n11408) );
  INV_X8 U10561 ( .A(n6422), .ZN(n6423) );
  NAND2_X4 U10562 ( .A1(n11987), .A2(n11986), .ZN(n12435) );
  NAND2_X4 U10563 ( .A1(n10549), .A2(n10548), .ZN(n10917) );
  NAND3_X2 U10564 ( .A1(n10512), .A2(n10511), .A3(net361984), .ZN(n10549) );
  OAI22_X4 U10565 ( .A1(n11379), .A2(net368462), .B1(n11453), .B2(net368195), 
        .ZN(n11445) );
  MUX2_X2 U10566 ( .A(n7301), .B(n7300), .S(net366979), .Z(n7302) );
  NAND2_X4 U10567 ( .A1(n11517), .A2(n11516), .ZN(n11675) );
  NAND3_X2 U10568 ( .A1(n5893), .A2(n11550), .A3(n5008), .ZN(n11580) );
  NAND2_X2 U10569 ( .A1(n12004), .A2(n5943), .ZN(n12079) );
  NAND3_X2 U10570 ( .A1(n12296), .A2(n12297), .A3(n12283), .ZN(n12298) );
  NAND3_X2 U10571 ( .A1(net369287), .A2(n11127), .A3(n11128), .ZN(net361404)
         );
  XNOR2_X2 U10572 ( .A(n10745), .B(n10827), .ZN(n10751) );
  INV_X1 U10573 ( .A(n11701), .ZN(n11578) );
  NAND3_X2 U10574 ( .A1(n12440), .A2(n12439), .A3(n12438), .ZN(n12441) );
  NAND2_X4 U10575 ( .A1(n11922), .A2(n11923), .ZN(n11925) );
  NAND2_X4 U10576 ( .A1(n11329), .A2(n11408), .ZN(n11839) );
  OAI21_X1 U10577 ( .B1(n5989), .B2(n6386), .A(n12357), .ZN(n12195) );
  INV_X8 U10578 ( .A(n11279), .ZN(n6424) );
  INV_X16 U10579 ( .A(n6424), .ZN(n6425) );
  NAND4_X4 U10580 ( .A1(n11340), .A2(net361053), .A3(n11367), .A4(n11341), 
        .ZN(n11353) );
  NAND2_X1 U10581 ( .A1(n11364), .A2(net360631), .ZN(net361009) );
  NAND2_X4 U10582 ( .A1(aluBoi_multBoi_temppp[44]), .A2(n11363), .ZN(net360631) );
  NAND3_X2 U10583 ( .A1(n10621), .A2(n10714), .A3(net361949), .ZN(n10750) );
  NAND3_X2 U10584 ( .A1(n11915), .A2(n11916), .A3(n11914), .ZN(n11945) );
  NAND3_X2 U10585 ( .A1(n11914), .A2(n11915), .A3(n11916), .ZN(n11902) );
  NAND2_X4 U10586 ( .A1(n11205), .A2(n11206), .ZN(n11079) );
  INV_X1 U10587 ( .A(n11685), .ZN(n11666) );
  NOR2_X4 U10588 ( .A1(n11568), .A2(n11567), .ZN(n11561) );
  NOR4_X4 U10589 ( .A1(n11549), .A2(n6092), .A3(n11660), .A4(n11560), .ZN(
        n11568) );
  NAND3_X2 U10590 ( .A1(n12087), .A2(n12034), .A3(n12033), .ZN(n12035) );
  INV_X32 U10591 ( .A(net369248), .ZN(net369242) );
  INV_X32 U10592 ( .A(net369248), .ZN(net369244) );
  INV_X32 U10593 ( .A(net369248), .ZN(net369246) );
  INV_X32 U10594 ( .A(net369240), .ZN(net369234) );
  INV_X32 U10595 ( .A(net369240), .ZN(net369236) );
  INV_X32 U10596 ( .A(net369224), .ZN(net369218) );
  INV_X32 U10597 ( .A(net369224), .ZN(net369220) );
  INV_X32 U10598 ( .A(net369224), .ZN(net369222) );
  INV_X32 U10599 ( .A(net369158), .ZN(net369224) );
  INV_X32 U10600 ( .A(net369216), .ZN(net369212) );
  INV_X32 U10601 ( .A(net369216), .ZN(net369214) );
  INV_X16 U10602 ( .A(net368903), .ZN(net369206) );
  XNOR2_X2 U10603 ( .A(n11782), .B(n11781), .ZN(n6430) );
  NAND3_X2 U10604 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n6431) );
  INV_X16 U10605 ( .A(net369139), .ZN(net369145) );
  INV_X8 U10606 ( .A(net369140), .ZN(net369148) );
  INV_X8 U10607 ( .A(net369140), .ZN(net369149) );
  INV_X16 U10608 ( .A(net369160), .ZN(net369154) );
  INV_X16 U10609 ( .A(net369142), .ZN(net369155) );
  INV_X16 U10610 ( .A(net369142), .ZN(net369156) );
  INV_X16 U10611 ( .A(n5763), .ZN(net369157) );
  INV_X16 U10612 ( .A(net369160), .ZN(net369161) );
  INV_X16 U10613 ( .A(net369160), .ZN(net369162) );
  INV_X16 U10614 ( .A(net369160), .ZN(net369163) );
  INV_X16 U10615 ( .A(net369160), .ZN(net369164) );
  INV_X16 U10616 ( .A(n5763), .ZN(net369166) );
  OAI21_X4 U10617 ( .B1(n8183), .B2(n8182), .A(n8181), .ZN(net369137) );
  NOR2_X4 U10618 ( .A1(net362342), .A2(n8180), .ZN(n8181) );
  AOI21_X2 U10619 ( .B1(n5880), .B2(n11871), .A(n5996), .ZN(n11872) );
  OAI21_X2 U10620 ( .B1(n5995), .B2(n11762), .A(n11875), .ZN(n11837) );
  XNOR2_X2 U10621 ( .A(n5958), .B(n11456), .ZN(n6432) );
  XNOR2_X2 U10622 ( .A(n11943), .B(net360235), .ZN(net359911) );
  NAND2_X1 U10623 ( .A1(n9988), .A2(n9992), .ZN(n6434) );
  NAND2_X1 U10624 ( .A1(n9988), .A2(n9992), .ZN(MoLanBoJ) );
  NAND2_X4 U10625 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  NOR2_X4 U10626 ( .A1(n12467), .A2(n12466), .ZN(n12472) );
  OAI21_X4 U10627 ( .B1(n11970), .B2(n12518), .A(net359905), .ZN(n11971) );
  OAI21_X2 U10628 ( .B1(n10701), .B2(net368467), .A(n10700), .ZN(n10702) );
  AND2_X2 U10629 ( .A1(net359809), .A2(net359495), .ZN(n6438) );
  NAND2_X4 U10630 ( .A1(n10454), .A2(n10453), .ZN(net362257) );
  NOR2_X2 U10631 ( .A1(n12542), .A2(n12541), .ZN(n12546) );
  NAND2_X4 U10632 ( .A1(n10728), .A2(n6440), .ZN(n10790) );
  INV_X4 U10633 ( .A(n6439), .ZN(n6440) );
  NAND2_X4 U10634 ( .A1(n10613), .A2(n10689), .ZN(n10633) );
  NAND2_X2 U10635 ( .A1(n6425), .A2(n11376), .ZN(n11224) );
  AOI22_X2 U10636 ( .A1(n11592), .A2(n11798), .B1(n11798), .B2(n5887), .ZN(
        n11622) );
  NAND2_X1 U10637 ( .A1(n10951), .A2(n10950), .ZN(net361417) );
  AOI21_X1 U10638 ( .B1(n9857), .B2(n9856), .A(n8031), .ZN(n7752) );
  INV_X8 U10639 ( .A(n8031), .ZN(n9855) );
  OAI21_X2 U10640 ( .B1(n12117), .B2(n12116), .A(n12127), .ZN(n12128) );
  INV_X2 U10641 ( .A(n12115), .ZN(n12116) );
  NAND2_X4 U10642 ( .A1(n6154), .A2(n12096), .ZN(n12127) );
  XNOR2_X2 U10643 ( .A(n10734), .B(n10733), .ZN(n6442) );
  NAND2_X4 U10644 ( .A1(n12383), .A2(n12382), .ZN(n12449) );
  INV_X2 U10645 ( .A(n12039), .ZN(n12051) );
  OAI22_X4 U10646 ( .A1(n11975), .A2(net368462), .B1(n12064), .B2(net368195), 
        .ZN(n11995) );
  NAND2_X4 U10647 ( .A1(n5151), .A2(n10914), .ZN(n10726) );
  NAND2_X4 U10648 ( .A1(n11697), .A2(net360583), .ZN(n12225) );
  NOR2_X1 U10649 ( .A1(net362287), .A2(n6574), .ZN(n10404) );
  AOI21_X1 U10650 ( .B1(n5288), .B2(net362287), .A(n5386), .ZN(n9682) );
  OAI21_X4 U10651 ( .B1(n12101), .B2(n4985), .A(n12418), .ZN(n12134) );
  XNOR2_X1 U10652 ( .A(n6565), .B(net362287), .ZN(n8711) );
  NAND2_X4 U10653 ( .A1(n11658), .A2(n11657), .ZN(n11849) );
  NOR2_X1 U10654 ( .A1(n11067), .A2(n6067), .ZN(n11069) );
  NAND2_X4 U10655 ( .A1(n11604), .A2(n11603), .ZN(n11827) );
  NAND2_X4 U10656 ( .A1(n11755), .A2(net360513), .ZN(n11875) );
  NAND2_X2 U10657 ( .A1(n12038), .A2(n12381), .ZN(n12083) );
  NAND2_X4 U10658 ( .A1(n12481), .A2(net129670), .ZN(n12548) );
  NAND3_X2 U10659 ( .A1(n11773), .A2(n11978), .A3(n11977), .ZN(n12055) );
  NAND2_X4 U10660 ( .A1(n9452), .A2(n9453), .ZN(n9751) );
  NAND3_X1 U10661 ( .A1(n12279), .A2(n12278), .A3(n12353), .ZN(n12370) );
  NAND2_X4 U10662 ( .A1(n12278), .A2(n12353), .ZN(n12189) );
  NAND3_X2 U10663 ( .A1(n11271), .A2(n11399), .A3(n11402), .ZN(n11208) );
  NAND2_X4 U10664 ( .A1(n12236), .A2(n12240), .ZN(n12448) );
  NAND2_X4 U10665 ( .A1(n11428), .A2(n11427), .ZN(n11495) );
  NOR3_X4 U10666 ( .A1(n11403), .A2(n6425), .A3(n6422), .ZN(n11280) );
  NAND3_X2 U10667 ( .A1(net361829), .A2(n10855), .A3(net361828), .ZN(n10798)
         );
  OAI21_X2 U10668 ( .B1(net361748), .B2(net376691), .A(n10855), .ZN(n10799) );
  NAND2_X4 U10669 ( .A1(net361889), .A2(net361536), .ZN(net361835) );
  NAND2_X4 U10670 ( .A1(n12538), .A2(n5988), .ZN(net359470) );
  INV_X2 U10671 ( .A(n12538), .ZN(n12539) );
  NAND3_X2 U10672 ( .A1(n11414), .A2(n11410), .A3(n11409), .ZN(n11334) );
  OAI211_X4 U10673 ( .C1(n12050), .C2(n12051), .A(n12049), .B(n12174), .ZN(
        n12255) );
  NOR2_X2 U10674 ( .A1(n12100), .A2(n12030), .ZN(n12036) );
  NAND2_X4 U10675 ( .A1(n11538), .A2(n11542), .ZN(n11539) );
  NAND2_X1 U10676 ( .A1(n10905), .A2(n11229), .ZN(n10743) );
  NAND3_X2 U10677 ( .A1(n11232), .A2(n10906), .A3(n10905), .ZN(n10907) );
  NAND2_X4 U10678 ( .A1(n12386), .A2(n12282), .ZN(n12394) );
  OAI22_X4 U10679 ( .A1(n5305), .A2(net368462), .B1(n6076), .B2(net368195), 
        .ZN(n11620) );
  INV_X8 U10680 ( .A(n11094), .ZN(n10947) );
  NAND2_X4 U10681 ( .A1(net362239), .A2(net377611), .ZN(n10578) );
  AOI21_X2 U10682 ( .B1(n12113), .B2(n6048), .A(n12111), .ZN(n12129) );
  INV_X2 U10683 ( .A(n9097), .ZN(n9098) );
  XNOR2_X1 U10684 ( .A(n9751), .B(n9750), .ZN(n9753) );
  NAND2_X4 U10685 ( .A1(n9750), .A2(n9751), .ZN(n9741) );
  NAND2_X4 U10686 ( .A1(n9094), .A2(n9097), .ZN(n9101) );
  INV_X2 U10687 ( .A(n12393), .ZN(n12395) );
  NAND3_X2 U10688 ( .A1(n11059), .A2(n10727), .A3(n11192), .ZN(n10791) );
  NAND3_X2 U10689 ( .A1(n11059), .A2(n11192), .A3(n10727), .ZN(n11000) );
  NAND2_X4 U10690 ( .A1(n12245), .A2(n6033), .ZN(n12284) );
  NAND2_X4 U10691 ( .A1(n12115), .A2(n12114), .ZN(n12245) );
  NAND2_X1 U10692 ( .A1(n10771), .A2(n10770), .ZN(n10772) );
  OAI21_X1 U10693 ( .B1(n6562), .B2(n9626), .A(n10724), .ZN(n9630) );
  OAI21_X1 U10694 ( .B1(n5007), .B2(n6563), .A(n6560), .ZN(n9627) );
  NAND2_X1 U10695 ( .A1(n8588), .A2(n10724), .ZN(n9075) );
  INV_X1 U10696 ( .A(n13525), .ZN(n10500) );
  INV_X1 U10697 ( .A(n13525), .ZN(n10581) );
  INV_X1 U10698 ( .A(n10579), .ZN(n10499) );
  INV_X8 U10699 ( .A(n6414), .ZN(n6798) );
  NOR3_X2 U10700 ( .A1(net362256), .A2(n10461), .A3(net362224), .ZN(n10463) );
  NAND2_X2 U10701 ( .A1(n12391), .A2(n12160), .ZN(n12534) );
  NOR2_X1 U10702 ( .A1(n11689), .A2(n6082), .ZN(n11690) );
  INV_X8 U10703 ( .A(n12235), .ZN(n12451) );
  NAND2_X4 U10704 ( .A1(n10838), .A2(net378405), .ZN(n10824) );
  OAI211_X4 U10705 ( .C1(n11911), .C2(n12090), .A(n12107), .B(n12089), .ZN(
        n12145) );
  NAND2_X4 U10706 ( .A1(n11463), .A2(n11462), .ZN(n11613) );
  NOR2_X2 U10707 ( .A1(n6251), .A2(n10573), .ZN(n10458) );
  INV_X4 U10708 ( .A(n12548), .ZN(n12549) );
  INV_X2 U10709 ( .A(n12369), .ZN(n12280) );
  NAND2_X1 U10710 ( .A1(n6095), .A2(n11641), .ZN(n11387) );
  NAND3_X2 U10711 ( .A1(n11400), .A2(n11458), .A3(n11641), .ZN(n11405) );
  NAND3_X2 U10712 ( .A1(n11646), .A2(n11593), .A3(n11374), .ZN(n11629) );
  NAND3_X2 U10713 ( .A1(n11578), .A2(n11703), .A3(n11850), .ZN(n11869) );
  NAND2_X4 U10714 ( .A1(n12419), .A2(n12418), .ZN(n12391) );
  NAND2_X1 U10715 ( .A1(n5965), .A2(n11024), .ZN(n10796) );
  NAND2_X4 U10716 ( .A1(n8700), .A2(net362253), .ZN(n10579) );
  NAND2_X4 U10717 ( .A1(n11839), .A2(n11409), .ZN(n11346) );
  NAND2_X4 U10718 ( .A1(n9469), .A2(n9470), .ZN(n8883) );
  NAND2_X4 U10719 ( .A1(n11550), .A2(n5964), .ZN(n11538) );
  INV_X8 U10720 ( .A(n11659), .ZN(n11855) );
  NAND2_X4 U10721 ( .A1(n8880), .A2(n9080), .ZN(n9087) );
  OAI21_X2 U10722 ( .B1(net359809), .B2(net359495), .A(net100619), .ZN(n12308)
         );
  NAND2_X4 U10723 ( .A1(n10624), .A2(n10617), .ZN(n10714) );
  NAND3_X4 U10724 ( .A1(n11206), .A2(n11205), .A3(n11204), .ZN(n11409) );
  NAND2_X4 U10725 ( .A1(n11077), .A2(n6425), .ZN(n11205) );
  OAI211_X4 U10726 ( .C1(n11969), .C2(n11968), .A(n11967), .B(
        aluBoi_multBoi_temppp[55]), .ZN(net359905) );
  INV_X8 U10727 ( .A(n10974), .ZN(n10980) );
  NAND2_X4 U10728 ( .A1(n12505), .A2(n12506), .ZN(n12504) );
  NAND2_X4 U10729 ( .A1(net361032), .A2(net361033), .ZN(net361002) );
  INV_X2 U10730 ( .A(net361021), .ZN(net361032) );
  INV_X8 U10731 ( .A(n11840), .ZN(n11842) );
  NAND3_X4 U10732 ( .A1(n11353), .A2(n11352), .A3(n11365), .ZN(n11348) );
  NAND2_X4 U10733 ( .A1(n11507), .A2(n11560), .ZN(n11564) );
  NAND3_X2 U10734 ( .A1(net362240), .A2(net362178), .A3(net361984), .ZN(n10502) );
  NOR2_X4 U10735 ( .A1(n11713), .A2(n6277), .ZN(n11406) );
  NAND3_X4 U10736 ( .A1(n11106), .A2(n11105), .A3(n5121), .ZN(n11154) );
  INV_X8 U10737 ( .A(n10617), .ZN(n10627) );
  NAND2_X4 U10738 ( .A1(n10729), .A2(n11230), .ZN(n10949) );
  NAND2_X4 U10739 ( .A1(n10712), .A2(n10713), .ZN(n10827) );
  NAND3_X2 U10740 ( .A1(n11906), .A2(n11904), .A3(n11905), .ZN(n12108) );
  NAND4_X4 U10741 ( .A1(n10570), .A2(net362287), .A3(n10520), .A4(net362224), 
        .ZN(net362239) );
  NAND2_X4 U10742 ( .A1(net361022), .A2(net361031), .ZN(n11350) );
  NAND2_X4 U10743 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  NAND2_X2 U10744 ( .A1(net360017), .A2(n12132), .ZN(n12531) );
  NAND2_X4 U10745 ( .A1(n12194), .A2(n11988), .ZN(n12028) );
  NAND2_X4 U10746 ( .A1(n12107), .A2(n12127), .ZN(n12100) );
  NAND2_X4 U10747 ( .A1(n11783), .A2(n11800), .ZN(n11788) );
  NAND2_X4 U10748 ( .A1(n11779), .A2(n6216), .ZN(n11783) );
  NAND2_X1 U10749 ( .A1(net359524), .A2(net100619), .ZN(n12516) );
  NAND2_X4 U10750 ( .A1(net359524), .A2(net360011), .ZN(n12519) );
  OAI211_X1 U10751 ( .C1(net361318), .C2(net361319), .A(
        aluBoi_multBoi_temppp[41]), .B(net361320), .ZN(net359788) );
  NAND3_X2 U10752 ( .A1(net377501), .A2(n11163), .A3(n5047), .ZN(net361276) );
  NAND2_X4 U10753 ( .A1(net361814), .A2(n5769), .ZN(n10762) );
  NAND3_X2 U10754 ( .A1(n11696), .A2(aluBoi_multBoi_temppp[51]), .A3(n5080), 
        .ZN(net359535) );
  NAND2_X2 U10755 ( .A1(n11696), .A2(n11940), .ZN(n11937) );
  NAND2_X1 U10756 ( .A1(n11690), .A2(n11960), .ZN(n11694) );
  NAND3_X2 U10757 ( .A1(n11860), .A2(n11861), .A3(n11862), .ZN(n11865) );
  NAND2_X4 U10758 ( .A1(n9735), .A2(n9736), .ZN(n9452) );
  AOI22_X4 U10759 ( .A1(n9044), .A2(n9045), .B1(n9009), .B2(n6521), .ZN(n9116)
         );
  NAND2_X1 U10760 ( .A1(n9102), .A2(n9100), .ZN(n9073) );
  OAI211_X4 U10761 ( .C1(n12091), .C2(n12090), .A(n12089), .B(n12088), .ZN(
        n12133) );
  OAI21_X2 U10762 ( .B1(n11898), .B2(n11897), .A(n11896), .ZN(n11916) );
  NOR2_X1 U10763 ( .A1(n11896), .A2(n11897), .ZN(n11894) );
  NAND2_X4 U10764 ( .A1(n11275), .A2(n11274), .ZN(n11420) );
  NAND2_X4 U10765 ( .A1(n11836), .A2(n11955), .ZN(n12094) );
  OAI21_X2 U10766 ( .B1(n11359), .B2(n11358), .A(n11357), .ZN(net361020) );
  INV_X2 U10767 ( .A(net362159), .ZN(net362156) );
  NOR2_X4 U10768 ( .A1(n12549), .A2(net359451), .ZN(n12554) );
  NAND2_X4 U10769 ( .A1(n6129), .A2(n11586), .ZN(n11797) );
  NAND2_X4 U10770 ( .A1(n12232), .A2(n12233), .ZN(n12241) );
  OAI21_X4 U10771 ( .B1(n12194), .B2(n12193), .A(n12192), .ZN(n12369) );
  NAND2_X4 U10772 ( .A1(n11226), .A2(n11225), .ZN(n11375) );
  NAND2_X2 U10773 ( .A1(n7150), .A2(net367025), .ZN(n6499) );
  NAND2_X1 U10774 ( .A1(n11036), .A2(n10989), .ZN(n10938) );
  NAND2_X1 U10775 ( .A1(n10772), .A2(n5947), .ZN(n10853) );
  AOI22_X1 U10776 ( .A1(n9731), .A2(aluBoi_aluBoi_shft_sraout[31]), .B1(n5766), 
        .B2(n9779), .ZN(n9783) );
  XNOR2_X1 U10777 ( .A(n9781), .B(n5766), .ZN(n9782) );
  XNOR2_X1 U10778 ( .A(n5978), .B(n9115), .ZN(n13140) );
  NAND2_X4 U10779 ( .A1(n6034), .A2(n12291), .ZN(n12418) );
  INV_X8 U10780 ( .A(n12030), .ZN(n12292) );
  OAI211_X4 U10781 ( .C1(n7806), .C2(n7805), .A(net361491), .B(n7804), .ZN(
        n10704) );
  NAND4_X4 U10782 ( .A1(n11705), .A2(n11703), .A3(n11704), .A4(n11856), .ZN(
        n11840) );
  NAND2_X4 U10783 ( .A1(n10890), .A2(n10722), .ZN(n11249) );
  NAND2_X4 U10784 ( .A1(n5935), .A2(n5939), .ZN(n11282) );
  NAND2_X4 U10785 ( .A1(n11829), .A2(n12039), .ZN(n12069) );
  NAND2_X2 U10786 ( .A1(n12543), .A2(net359418), .ZN(n12551) );
  NAND3_X2 U10787 ( .A1(net362297), .A2(n7638), .A3(n7637), .ZN(n7639) );
  OAI22_X4 U10788 ( .A1(net360723), .A2(net368462), .B1(net368195), .B2(
        net360403), .ZN(n11717) );
  NAND2_X4 U10789 ( .A1(n6012), .A2(n11606), .ZN(net360403) );
  NAND2_X4 U10790 ( .A1(n12263), .A2(n12264), .ZN(n12353) );
  NAND3_X4 U10791 ( .A1(n11527), .A2(n11528), .A3(n11609), .ZN(n11530) );
  NAND3_X1 U10792 ( .A1(net359533), .A2(n12510), .A3(net377689), .ZN(n12512)
         );
  NOR2_X1 U10793 ( .A1(n11319), .A2(n5942), .ZN(n11165) );
  NAND3_X2 U10794 ( .A1(net361899), .A2(net361835), .A3(net361886), .ZN(
        net361357) );
  NAND2_X4 U10795 ( .A1(n10569), .A2(n10722), .ZN(n11301) );
  OAI22_X4 U10796 ( .A1(n12138), .A2(n12137), .B1(n12136), .B2(n12135), .ZN(
        net360033) );
  NAND2_X4 U10797 ( .A1(n6070), .A2(net129670), .ZN(n12538) );
  NAND2_X4 U10798 ( .A1(net362256), .A2(net362224), .ZN(n10573) );
  NAND2_X4 U10799 ( .A1(n12158), .A2(n12157), .ZN(n12408) );
  XNOR2_X1 U10800 ( .A(n9092), .B(n9091), .ZN(n12973) );
  NAND2_X1 U10801 ( .A1(n9741), .A2(n9740), .ZN(n9762) );
  NAND2_X4 U10802 ( .A1(n9091), .A2(n8718), .ZN(n9093) );
  INV_X8 U10803 ( .A(net360927), .ZN(net360617) );
  NAND2_X4 U10804 ( .A1(aluBoi_multBoi_temppp[59]), .A2(n12084), .ZN(net359501) );
  NAND2_X1 U10805 ( .A1(n12093), .A2(n12086), .ZN(n11911) );
  NAND2_X1 U10806 ( .A1(n12086), .A2(n12093), .ZN(n12091) );
  NAND2_X4 U10807 ( .A1(n10833), .A2(n10834), .ZN(n10958) );
  NAND3_X1 U10808 ( .A1(n5937), .A2(n6004), .A3(n12449), .ZN(n12410) );
  NOR2_X1 U10809 ( .A1(net377453), .A2(net359531), .ZN(n12511) );
  NAND3_X1 U10810 ( .A1(n5080), .A2(n5975), .A3(aluBoi_multBoi_temppp[52]), 
        .ZN(n11939) );
  NAND2_X4 U10811 ( .A1(n11548), .A2(n11547), .ZN(n11862) );
  NAND3_X2 U10812 ( .A1(n11035), .A2(n6029), .A3(n5882), .ZN(n11092) );
  XNOR2_X1 U10813 ( .A(n13525), .B(n9677), .ZN(n8702) );
  NAND2_X1 U10814 ( .A1(net360904), .A2(n10579), .ZN(n10533) );
  NAND2_X4 U10815 ( .A1(net360002), .A2(n12152), .ZN(n12205) );
  NAND2_X4 U10816 ( .A1(n11548), .A2(n11839), .ZN(n11699) );
  NAND2_X4 U10817 ( .A1(n11709), .A2(n11389), .ZN(n11624) );
  NAND3_X4 U10818 ( .A1(n11050), .A2(n6061), .A3(n11049), .ZN(n11709) );
  NAND2_X4 U10819 ( .A1(n11193), .A2(n11192), .ZN(n10912) );
  XNOR2_X1 U10820 ( .A(n13219), .B(n5927), .ZN(n9457) );
  NOR2_X1 U10821 ( .A1(n5392), .A2(n13222), .ZN(n9733) );
  INV_X2 U10822 ( .A(n9093), .ZN(n9096) );
  XOR2_X1 U10823 ( .A(n9768), .B(n9767), .Z(n9771) );
  NAND3_X1 U10824 ( .A1(n9102), .A2(n9101), .A3(n9100), .ZN(n9106) );
  NAND2_X1 U10825 ( .A1(n9101), .A2(n9072), .ZN(n9074) );
  NAND2_X1 U10826 ( .A1(n9101), .A2(n9075), .ZN(n9066) );
  NAND2_X4 U10827 ( .A1(aluBoi_multBoi_temppp[56]), .A2(n12139), .ZN(net359486) );
  NAND2_X4 U10828 ( .A1(n10719), .A2(n10720), .ZN(n10745) );
  OAI211_X4 U10829 ( .C1(n11406), .C2(n11405), .A(n11640), .B(n11404), .ZN(
        n11500) );
  NAND4_X1 U10830 ( .A1(n11956), .A2(n12033), .A3(n11955), .A4(n12031), .ZN(
        n11957) );
  NAND3_X1 U10831 ( .A1(n11007), .A2(n6150), .A3(n5438), .ZN(n11018) );
  NAND3_X1 U10832 ( .A1(n5438), .A2(n11010), .A3(n6150), .ZN(n11016) );
  NAND3_X1 U10833 ( .A1(n6150), .A2(n11049), .A3(n11010), .ZN(n10992) );
  NAND3_X1 U10834 ( .A1(n11059), .A2(n11192), .A3(net368201), .ZN(n11195) );
  NAND2_X4 U10835 ( .A1(n11398), .A2(n11397), .ZN(n11459) );
  INV_X8 U10836 ( .A(n11043), .ZN(n11398) );
  NAND2_X4 U10837 ( .A1(n11879), .A2(n11844), .ZN(n12014) );
  OAI211_X4 U10838 ( .C1(n5999), .C2(n11843), .A(n11842), .B(n11841), .ZN(
        n11879) );
  NAND2_X4 U10839 ( .A1(n10905), .A2(n10610), .ZN(n11071) );
  NAND3_X2 U10840 ( .A1(n9065), .A2(n8726), .A3(n9064), .ZN(n8725) );
  AOI22_X4 U10841 ( .A1(n9199), .A2(n9200), .B1(n9151), .B2(net368572), .ZN(
        n9380) );
  NAND2_X4 U10842 ( .A1(n11332), .A2(n11345), .ZN(net361022) );
  NAND2_X4 U10843 ( .A1(n10582), .A2(net362161), .ZN(n10837) );
  NAND4_X4 U10844 ( .A1(n10837), .A2(n10838), .A3(n10958), .A4(n10839), .ZN(
        n10970) );
  OAI221_X4 U10845 ( .B1(n12128), .B2(n12129), .C1(n12294), .C2(n12293), .A(
        n12284), .ZN(n12140) );
  NAND2_X1 U10846 ( .A1(net376321), .A2(net359676), .ZN(n12399) );
  NAND3_X2 U10847 ( .A1(n11661), .A2(n11862), .A3(n11861), .ZN(n11895) );
  NOR2_X1 U10848 ( .A1(n11740), .A2(n11735), .ZN(n11259) );
  NAND2_X4 U10849 ( .A1(n11862), .A2(n11861), .ZN(n11549) );
  NAND2_X1 U10850 ( .A1(net368215), .A2(n6194), .ZN(n10705) );
  INV_X2 U10851 ( .A(net368926), .ZN(net368927) );
  INV_X16 U10852 ( .A(n13707), .ZN(n6508) );
  INV_X2 U10853 ( .A(n6444), .ZN(n6445) );
  NAND2_X1 U10854 ( .A1(regBoiz_regfile_25__9_), .A2(n6736), .ZN(n541) );
  NAND2_X1 U10855 ( .A1(regBoiz_regfile_28__9_), .A2(n6748), .ZN(n440) );
  INV_X2 U10856 ( .A(n6446), .ZN(n6447) );
  NAND2_X4 U10857 ( .A1(net361491), .A2(n7183), .ZN(n11771) );
  NAND2_X1 U10858 ( .A1(regBoiz_regfile_28__4_), .A2(n6747), .ZN(n445) );
  NAND2_X1 U10859 ( .A1(regBoiz_regfile_13__4_), .A2(n6690), .ZN(n981) );
  MUX2_X1 U10860 ( .A(regBoiz_regfile_10__4_), .B(regBoiz_regfile_11__4_), .S(
        net369165), .Z(n9315) );
  INV_X2 U10861 ( .A(n6448), .ZN(n6449) );
  INV_X2 U10862 ( .A(n6450), .ZN(n6451) );
  INV_X2 U10863 ( .A(n6452), .ZN(n6453) );
  MUX2_X1 U10864 ( .A(regBoiz_regfile_14__4_), .B(regBoiz_regfile_15__4_), .S(
        net369162), .Z(n9317) );
  NAND2_X1 U10865 ( .A1(regBoiz_regfile_14__4_), .A2(n6695), .ZN(n948) );
  NAND2_X1 U10866 ( .A1(regBoiz_regfile_25__4_), .A2(n6738), .ZN(n546) );
  MUX2_X1 U10867 ( .A(regBoiz_regfile_26__4_), .B(regBoiz_regfile_27__4_), .S(
        net369166), .Z(n9329) );
  NAND2_X1 U10868 ( .A1(regBoiz_regfile_26__4_), .A2(n6742), .ZN(n513) );
  INV_X2 U10869 ( .A(n6455), .ZN(n6456) );
  OAI21_X2 U10870 ( .B1(n6659), .B2(n6748), .A(n440), .ZN(n3791) );
  OAI21_X2 U10871 ( .B1(n6669), .B2(n6747), .A(n445), .ZN(n3626) );
  INV_X8 U10872 ( .A(net368712), .ZN(net368713) );
  NAND2_X1 U10873 ( .A1(regBoiz_regfile_15__10_), .A2(n6699), .ZN(n939) );
  MUX2_X1 U10874 ( .A(n7773), .B(n7772), .S(net366973), .Z(n7774) );
  MUX2_X2 U10875 ( .A(n7253), .B(n7254), .S(net368862), .Z(n7258) );
  NAND2_X1 U10876 ( .A1(regBoiz_regfile_15__7_), .A2(n6697), .ZN(n911) );
  NAND2_X1 U10877 ( .A1(regBoiz_regfile_29__10_), .A2(n6751), .ZN(n437) );
  INV_X4 U10878 ( .A(n6477), .ZN(n7263) );
  INV_X4 U10879 ( .A(n6483), .ZN(n7267) );
  INV_X4 U10880 ( .A(n6495), .ZN(n7085) );
  NAND2_X1 U10881 ( .A1(regBoiz_regfile_27__10_), .A2(n6745), .ZN(n504) );
  NAND2_X1 U10882 ( .A1(regBoiz_regfile_23__10_), .A2(n6730), .ZN(n639) );
  MUX2_X2 U10883 ( .A(n6458), .B(n6459), .S(net367035), .Z(n6457) );
  INV_X2 U10884 ( .A(n6460), .ZN(n6461) );
  NAND3_X1 U10885 ( .A1(net362387), .A2(n8074), .A3(n8049), .ZN(n8057) );
  NOR2_X1 U10886 ( .A1(n8074), .A2(n5510), .ZN(n8088) );
  INV_X2 U10887 ( .A(n6463), .ZN(n6464) );
  INV_X4 U10888 ( .A(n6470), .ZN(n7300) );
  INV_X2 U10889 ( .A(n6465), .ZN(n6466) );
  INV_X2 U10890 ( .A(n6467), .ZN(n6468) );
  MUX2_X2 U10891 ( .A(n6471), .B(n6472), .S(net367035), .Z(n6470) );
  INV_X16 U10892 ( .A(net368713), .ZN(net367039) );
  NAND2_X1 U10893 ( .A1(regBoiz_regfile_31__10_), .A2(n6757), .ZN(n337) );
  OAI211_X4 U10894 ( .C1(n7348), .C2(n7347), .A(net361491), .B(n7346), .ZN(
        n9813) );
  NAND2_X1 U10895 ( .A1(n7210), .A2(net376063), .ZN(n6474) );
  NAND2_X2 U10896 ( .A1(n6473), .A2(n6474), .ZN(n7212) );
  NAND2_X4 U10897 ( .A1(n6998), .A2(n6997), .ZN(net364882) );
  INV_X8 U10898 ( .A(net364882), .ZN(net365336) );
  NAND2_X4 U10899 ( .A1(net364968), .A2(daddr[3]), .ZN(net362253) );
  INV_X8 U10900 ( .A(n9893), .ZN(n11243) );
  MUX2_X1 U10901 ( .A(n7374), .B(n7373), .S(net366927), .Z(n7375) );
  MUX2_X1 U10902 ( .A(n7404), .B(n7403), .S(net366927), .Z(n7405) );
  INV_X4 U10903 ( .A(n6500), .ZN(n7269) );
  AOI22_X2 U10904 ( .A1(regBoiz_regfile_9__12_), .A2(net367003), .B1(
        regBoiz_regfile_11__12_), .B2(net366985), .ZN(n7355) );
  NAND2_X1 U10905 ( .A1(regBoiz_regfile_17__12_), .A2(net367001), .ZN(n6475)
         );
  NAND2_X1 U10906 ( .A1(regBoiz_regfile_19__12_), .A2(net366985), .ZN(n6476)
         );
  AND2_X2 U10907 ( .A1(n6475), .A2(n6476), .ZN(n7363) );
  OAI22_X1 U10908 ( .A1(n7364), .A2(net375713), .B1(n7363), .B2(net367043), 
        .ZN(n7368) );
  OAI22_X1 U10909 ( .A1(n7352), .A2(net367031), .B1(n7351), .B2(net367043), 
        .ZN(n7353) );
  AOI22_X2 U10910 ( .A1(regBoiz_regfile_5__12_), .A2(net367003), .B1(
        regBoiz_regfile_7__12_), .B2(net366985), .ZN(n7351) );
  AOI22_X1 U10911 ( .A1(regBoiz_regfile_0__13_), .A2(net367001), .B1(
        regBoiz_regfile_2__13_), .B2(net366985), .ZN(n7381) );
  AOI22_X1 U10912 ( .A1(regBoiz_regfile_0__12_), .A2(net367003), .B1(
        regBoiz_regfile_2__12_), .B2(net366985), .ZN(n7350) );
  AOI22_X1 U10913 ( .A1(regBoiz_regfile_1__13_), .A2(net367003), .B1(
        regBoiz_regfile_3__13_), .B2(net366985), .ZN(n7380) );
  AOI22_X1 U10914 ( .A1(regBoiz_regfile_16__12_), .A2(net367003), .B1(
        regBoiz_regfile_18__12_), .B2(net366985), .ZN(n7364) );
  AOI22_X1 U10915 ( .A1(regBoiz_regfile_0__29_), .A2(net366907), .B1(
        regBoiz_regfile_8__29_), .B2(net377464), .ZN(n8051) );
  MUX2_X2 U10916 ( .A(n6478), .B(n6479), .S(net376574), .Z(n6477) );
  MUX2_X2 U10917 ( .A(n6481), .B(n6482), .S(net366901), .Z(n6480) );
  MUX2_X2 U10918 ( .A(n7270), .B(n7269), .S(net366981), .Z(n7271) );
  MUX2_X2 U10919 ( .A(n6484), .B(n6485), .S(net376541), .Z(n6483) );
  MUX2_X2 U10920 ( .A(n6487), .B(n6488), .S(net366907), .Z(n6486) );
  MUX2_X2 U10921 ( .A(n6490), .B(n6491), .S(net366905), .Z(n6489) );
  NAND2_X4 U10922 ( .A1(n9896), .A2(n6536), .ZN(n9897) );
  NAND2_X2 U10923 ( .A1(n7182), .A2(n6492), .ZN(n6493) );
  NAND2_X2 U10924 ( .A1(n7181), .A2(n6785), .ZN(n6494) );
  MUX2_X2 U10925 ( .A(n6496), .B(n6497), .S(net375929), .Z(n6495) );
  NAND2_X1 U10926 ( .A1(net363049), .A2(net368548), .ZN(n9876) );
  NAND2_X4 U10927 ( .A1(net361491), .A2(n7409), .ZN(n9842) );
  INV_X16 U10928 ( .A(n9898), .ZN(n11609) );
  NAND2_X2 U10929 ( .A1(n7151), .A2(net375614), .ZN(n6498) );
  NAND2_X2 U10930 ( .A1(n6499), .A2(n6498), .ZN(n7152) );
  MUX2_X2 U10931 ( .A(n6501), .B(n6502), .S(net375929), .Z(n6500) );
  MUX2_X2 U10932 ( .A(n6504), .B(n6505), .S(net376642), .Z(n6503) );
  NAND2_X4 U10933 ( .A1(n10570), .A2(n9785), .ZN(n11303) );
  NOR3_X2 U10934 ( .A1(n9784), .A2(net368498), .A3(net362362), .ZN(n9785) );
  INV_X8 U10935 ( .A(n8074), .ZN(n8157) );
  NAND2_X4 U10936 ( .A1(net365335), .A2(net365336), .ZN(n8074) );
  NAND2_X4 U10937 ( .A1(net361491), .A2(n7093), .ZN(n9802) );
  INV_X4 U10938 ( .A(net369316), .ZN(net367045) );
  NOR3_X1 U10939 ( .A1(n6194), .A2(n11194), .A3(net368209), .ZN(n11060) );
  INV_X8 U10940 ( .A(n11194), .ZN(n11232) );
  INV_X2 U10941 ( .A(net362253), .ZN(net362251) );
  NAND3_X1 U10942 ( .A1(n10479), .A2(n10478), .A3(net362253), .ZN(n10480) );
  NAND3_X1 U10943 ( .A1(n8103), .A2(net364905), .A3(net364904), .ZN(net364871)
         );
  NAND2_X4 U10944 ( .A1(n7152), .A2(net361491), .ZN(n9798) );
  INV_X16 U10945 ( .A(net368713), .ZN(net367035) );
  NAND2_X4 U10946 ( .A1(n7308), .A2(net361491), .ZN(n11520) );
  INV_X8 U10947 ( .A(n13522), .ZN(n6528) );
  NOR2_X1 U10948 ( .A1(net366965), .A2(n5961), .ZN(n7686) );
  NOR2_X1 U10949 ( .A1(net366999), .A2(n5961), .ZN(n7693) );
  INV_X2 U10950 ( .A(n5960), .ZN(n8012) );
  INV_X2 U10951 ( .A(n5961), .ZN(n8015) );
  INV_X8 U10952 ( .A(n9880), .ZN(n7557) );
  INV_X8 U10953 ( .A(n11721), .ZN(n11304) );
  NAND2_X4 U10954 ( .A1(n11304), .A2(n11305), .ZN(n9898) );
  NAND2_X1 U10955 ( .A1(n10473), .A2(n6251), .ZN(n10586) );
  NAND2_X1 U10956 ( .A1(net345751), .A2(n6251), .ZN(n10544) );
  NAND2_X4 U10957 ( .A1(n12182), .A2(n12183), .ZN(n9903) );
  INV_X16 U10958 ( .A(net362175), .ZN(net361984) );
  NAND2_X4 U10959 ( .A1(net362253), .A2(net362265), .ZN(net362175) );
  NAND3_X2 U10960 ( .A1(net368571), .A2(n5305), .A3(n11718), .ZN(n9796) );
  NAND2_X1 U10961 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NAND3_X1 U10962 ( .A1(n11521), .A2(n11527), .A3(n11609), .ZN(n11522) );
  INV_X8 U10963 ( .A(MoLanBoJ), .ZN(n6548) );
  NAND2_X4 U10964 ( .A1(n7277), .A2(net361491), .ZN(n11720) );
  NAND2_X4 U10965 ( .A1(n7214), .A2(net361491), .ZN(n11727) );
  NAND2_X4 U10966 ( .A1(n9903), .A2(idOut_32_), .ZN(n9941) );
  INV_X32 U10967 ( .A(n6512), .ZN(n6513) );
  INV_X32 U10968 ( .A(n6516), .ZN(n6517) );
  INV_X32 U10969 ( .A(n13528), .ZN(n6520) );
  INV_X32 U10970 ( .A(n6520), .ZN(n6521) );
  NAND2_X4 U10971 ( .A1(n9813), .A2(n9815), .ZN(n13528) );
  INV_X32 U10972 ( .A(n6522), .ZN(n6523) );
  INV_X32 U10973 ( .A(n6524), .ZN(n6525) );
  NAND2_X4 U10974 ( .A1(n9843), .A2(n9844), .ZN(n13521) );
  INV_X32 U10975 ( .A(n6528), .ZN(n6529) );
  NAND2_X4 U10976 ( .A1(n7565), .A2(n9833), .ZN(n13533) );
  NAND2_X4 U10977 ( .A1(n7597), .A2(n9834), .ZN(n13531) );
  INV_X32 U10978 ( .A(n6538), .ZN(n6539) );
  NAND2_X4 U10979 ( .A1(n9895), .A2(n9894), .ZN(n13529) );
  INV_X32 U10980 ( .A(n6540), .ZN(n6541) );
  INV_X32 U10981 ( .A(n6546), .ZN(n6547) );
  INV_X32 U10982 ( .A(n8708), .ZN(n9718) );
  NAND2_X4 U10983 ( .A1(n5314), .A2(n5363), .ZN(n9677) );
  NAND2_X4 U10984 ( .A1(n10454), .A2(n10453), .ZN(n10560) );
  INV_X32 U10985 ( .A(n10139), .ZN(n10408) );
  INV_X32 U10986 ( .A(net368461), .ZN(net368462) );
  NAND2_X4 U10987 ( .A1(n5958), .A2(n5953), .ZN(n11400) );
  AND2_X4 U10988 ( .A1(n1209), .A2(n1147), .ZN(n1158) );
  INV_X32 U10989 ( .A(n6575), .ZN(n6573) );
  INV_X32 U10990 ( .A(n6575), .ZN(n6574) );
  INV_X16 U10991 ( .A(n10403), .ZN(n6575) );
  INV_X32 U10992 ( .A(net368213), .ZN(net368209) );
  INV_X32 U10993 ( .A(net368213), .ZN(net368211) );
  INV_X32 U10994 ( .A(net368217), .ZN(net368213) );
  INV_X32 U10995 ( .A(net368217), .ZN(net368215) );
  INV_X32 U10996 ( .A(net368201), .ZN(net368195) );
  INV_X32 U10997 ( .A(n6585), .ZN(n6581) );
  INV_X32 U10998 ( .A(n6585), .ZN(n6582) );
  INV_X32 U10999 ( .A(n6585), .ZN(n6583) );
  INV_X32 U11000 ( .A(n6585), .ZN(n6584) );
  INV_X32 U11001 ( .A(n6591), .ZN(n6589) );
  INV_X32 U11002 ( .A(n6586), .ZN(n6591) );
  INV_X32 U11003 ( .A(n6598), .ZN(n6595) );
  INV_X32 U11004 ( .A(n6599), .ZN(n6603) );
  INV_X32 U11005 ( .A(n6613), .ZN(n6612) );
  INV_X32 U11006 ( .A(n6617), .ZN(n6616) );
  INV_X32 U11007 ( .A(n6619), .ZN(n6618) );
  INV_X32 U11008 ( .A(net366995), .ZN(net366967) );
  INV_X32 U11009 ( .A(net366995), .ZN(net366969) );
  INV_X32 U11010 ( .A(net366991), .ZN(net366977) );
  INV_X32 U11011 ( .A(net366991), .ZN(net366979) );
  INV_X32 U11012 ( .A(net366991), .ZN(net366981) );
  INV_X32 U11013 ( .A(net367009), .ZN(net366995) );
  INV_X32 U11014 ( .A(net366947), .ZN(net366919) );
  INV_X32 U11015 ( .A(net366947), .ZN(net366921) );
  INV_X32 U11016 ( .A(net366945), .ZN(net366927) );
  INV_X32 U11017 ( .A(net366947), .ZN(net366933) );
  INV_X32 U11018 ( .A(net375310), .ZN(net366937) );
  INV_X32 U11019 ( .A(net366937), .ZN(net366945) );
  INV_X32 U11020 ( .A(n6790), .ZN(n6783) );
  INV_X32 U11021 ( .A(n6791), .ZN(n6784) );
  INV_X32 U11022 ( .A(n6791), .ZN(n6785) );
  INV_X32 U11023 ( .A(n6791), .ZN(n6786) );
  INV_X32 U11024 ( .A(n6790), .ZN(n6788) );
  INV_X32 U11025 ( .A(n6797), .ZN(n6791) );
  INV_X32 U11026 ( .A(n6817), .ZN(n6800) );
  INV_X32 U11027 ( .A(n6817), .ZN(n6801) );
  INV_X32 U11028 ( .A(n6817), .ZN(n6802) );
  INV_X32 U11029 ( .A(n6817), .ZN(n6804) );
  INV_X32 U11030 ( .A(n6814), .ZN(n6806) );
  INV_X32 U11031 ( .A(n6817), .ZN(n6807) );
  INV_X32 U11032 ( .A(n6817), .ZN(n6809) );
  INV_X32 U11033 ( .A(n6814), .ZN(n6810) );
  INV_X32 U11034 ( .A(n6814), .ZN(n6811) );
  INV_X32 U11035 ( .A(n6814), .ZN(n6812) );
  INV_X32 U11036 ( .A(n6814), .ZN(n6813) );
  INV_X32 U11037 ( .A(n6818), .ZN(n6817) );
  INV_X32 U11038 ( .A(n6827), .ZN(n6821) );
  INV_X32 U11039 ( .A(n6827), .ZN(n6822) );
  INV_X32 U11040 ( .A(n6824), .ZN(n6827) );
  INV_X32 U11041 ( .A(n5677), .ZN(n6830) );
  INV_X32 U11042 ( .A(n5344), .ZN(n6834) );
  NAND2_X2 U11043 ( .A1(didMult), .A2(n5691), .ZN(n9992) );
  NAND2_X2 U11044 ( .A1(n9992), .A2(n6959), .ZN(n13675) );
  NAND2_X2 U11045 ( .A1(n9992), .A2(n6943), .ZN(n13661) );
  MUX2_X2 U11046 ( .A(regBoiz_regfile_0__0_), .B(regBoiz_regfile_1__0_), .S(
        net367029), .Z(n6963) );
  MUX2_X2 U11047 ( .A(regBoiz_regfile_2__0_), .B(regBoiz_regfile_3__0_), .S(
        net376222), .Z(n6962) );
  MUX2_X2 U11048 ( .A(n6963), .B(n6962), .S(net366969), .Z(n6967) );
  MUX2_X2 U11049 ( .A(regBoiz_regfile_4__0_), .B(regBoiz_regfile_5__0_), .S(
        net367023), .Z(n6965) );
  MUX2_X2 U11050 ( .A(regBoiz_regfile_6__0_), .B(regBoiz_regfile_7__0_), .S(
        net367019), .Z(n6964) );
  MUX2_X2 U11051 ( .A(n6965), .B(n6964), .S(net366979), .Z(n6966) );
  MUX2_X2 U11052 ( .A(n6967), .B(n6966), .S(net366933), .Z(n6975) );
  MUX2_X2 U11053 ( .A(regBoiz_regfile_8__0_), .B(regBoiz_regfile_9__0_), .S(
        net367027), .Z(n6969) );
  MUX2_X2 U11054 ( .A(regBoiz_regfile_10__0_), .B(regBoiz_regfile_11__0_), .S(
        net375713), .Z(n6968) );
  MUX2_X2 U11055 ( .A(n6969), .B(n6968), .S(net366987), .Z(n6973) );
  MUX2_X2 U11056 ( .A(regBoiz_regfile_12__0_), .B(regBoiz_regfile_13__0_), .S(
        net375718), .Z(n6971) );
  MUX2_X2 U11057 ( .A(regBoiz_regfile_14__0_), .B(regBoiz_regfile_15__0_), .S(
        net367027), .Z(n6970) );
  MUX2_X2 U11058 ( .A(n6971), .B(n6970), .S(net366987), .Z(n6972) );
  MUX2_X2 U11059 ( .A(n6973), .B(n6972), .S(net366933), .Z(n6974) );
  MUX2_X2 U11060 ( .A(n6975), .B(n6974), .S(net375727), .Z(n6991) );
  MUX2_X2 U11061 ( .A(regBoiz_regfile_16__0_), .B(regBoiz_regfile_17__0_), .S(
        net367025), .Z(n6977) );
  MUX2_X2 U11062 ( .A(regBoiz_regfile_18__0_), .B(regBoiz_regfile_19__0_), .S(
        net367029), .Z(n6976) );
  MUX2_X2 U11063 ( .A(n6977), .B(n6976), .S(net366977), .Z(n6981) );
  MUX2_X2 U11064 ( .A(regBoiz_regfile_20__0_), .B(regBoiz_regfile_21__0_), .S(
        net367031), .Z(n6979) );
  MUX2_X2 U11065 ( .A(regBoiz_regfile_22__0_), .B(regBoiz_regfile_23__0_), .S(
        net367029), .Z(n6978) );
  MUX2_X2 U11066 ( .A(n6979), .B(n6978), .S(net366987), .Z(n6980) );
  MUX2_X2 U11067 ( .A(n6981), .B(n6980), .S(net366933), .Z(n6989) );
  MUX2_X2 U11068 ( .A(regBoiz_regfile_24__0_), .B(regBoiz_regfile_25__0_), .S(
        net375717), .Z(n6983) );
  MUX2_X2 U11069 ( .A(regBoiz_regfile_26__0_), .B(regBoiz_regfile_27__0_), .S(
        net367025), .Z(n6982) );
  MUX2_X2 U11070 ( .A(n6983), .B(n6982), .S(net366977), .Z(n6987) );
  MUX2_X2 U11071 ( .A(regBoiz_regfile_28__0_), .B(regBoiz_regfile_29__0_), .S(
        net367031), .Z(n6985) );
  MUX2_X2 U11072 ( .A(n6985), .B(n6984), .S(net366977), .Z(n6986) );
  MUX2_X2 U11073 ( .A(n6987), .B(n6986), .S(net366933), .Z(n6988) );
  MUX2_X2 U11074 ( .A(n6989), .B(n6988), .S(net369204), .Z(n6990) );
  MUX2_X2 U11075 ( .A(n6991), .B(n6990), .S(n5107), .Z(n6992) );
  INV_X4 U11076 ( .A(n6992), .ZN(n7000) );
  NOR2_X4 U11077 ( .A1(net366925), .A2(net369316), .ZN(n6993) );
  NOR2_X4 U11078 ( .A1(net369204), .A2(net366965), .ZN(n8144) );
  XNOR2_X2 U11079 ( .A(aluRw[2]), .B(net366927), .ZN(n6998) );
  NAND2_X2 U11080 ( .A1(net368221), .A2(daddr[31]), .ZN(n6999) );
  OAI21_X4 U11081 ( .B1(n7000), .B2(n5310), .A(n6999), .ZN(n13705) );
  MUX2_X2 U11082 ( .A(regBoiz_regfile_0__1_), .B(regBoiz_regfile_1__1_), .S(
        net367031), .Z(n7002) );
  MUX2_X2 U11083 ( .A(regBoiz_regfile_2__1_), .B(regBoiz_regfile_3__1_), .S(
        net375650), .Z(n7001) );
  MUX2_X2 U11084 ( .A(n7002), .B(n7001), .S(net366977), .Z(n7006) );
  MUX2_X2 U11085 ( .A(regBoiz_regfile_4__1_), .B(regBoiz_regfile_5__1_), .S(
        net375650), .Z(n7004) );
  MUX2_X2 U11086 ( .A(regBoiz_regfile_6__1_), .B(regBoiz_regfile_7__1_), .S(
        net367029), .Z(n7003) );
  MUX2_X2 U11087 ( .A(regBoiz_regfile_8__1_), .B(regBoiz_regfile_9__1_), .S(
        net367031), .Z(n7008) );
  MUX2_X2 U11088 ( .A(regBoiz_regfile_10__1_), .B(regBoiz_regfile_11__1_), .S(
        net375717), .Z(n7007) );
  MUX2_X2 U11089 ( .A(n7008), .B(n7007), .S(net366977), .Z(n7012) );
  MUX2_X2 U11090 ( .A(regBoiz_regfile_12__1_), .B(regBoiz_regfile_13__1_), .S(
        net376223), .Z(n7010) );
  MUX2_X2 U11091 ( .A(regBoiz_regfile_14__1_), .B(regBoiz_regfile_15__1_), .S(
        net376222), .Z(n7009) );
  MUX2_X2 U11092 ( .A(n7010), .B(n7009), .S(net366977), .Z(n7011) );
  MUX2_X2 U11093 ( .A(n7012), .B(n7011), .S(net366933), .Z(n7013) );
  MUX2_X2 U11094 ( .A(regBoiz_regfile_16__1_), .B(regBoiz_regfile_17__1_), .S(
        net367025), .Z(n7016) );
  MUX2_X2 U11095 ( .A(regBoiz_regfile_18__1_), .B(regBoiz_regfile_19__1_), .S(
        net367027), .Z(n7015) );
  MUX2_X2 U11096 ( .A(n7016), .B(n7015), .S(net366977), .Z(n7020) );
  MUX2_X2 U11097 ( .A(regBoiz_regfile_20__1_), .B(regBoiz_regfile_21__1_), .S(
        net367025), .Z(n7018) );
  MUX2_X2 U11098 ( .A(regBoiz_regfile_22__1_), .B(regBoiz_regfile_23__1_), .S(
        net367025), .Z(n7017) );
  MUX2_X2 U11099 ( .A(n7020), .B(n7019), .S(net366933), .Z(n7028) );
  MUX2_X2 U11100 ( .A(regBoiz_regfile_24__1_), .B(regBoiz_regfile_25__1_), .S(
        net367031), .Z(n7022) );
  MUX2_X2 U11101 ( .A(regBoiz_regfile_26__1_), .B(regBoiz_regfile_27__1_), .S(
        net367031), .Z(n7021) );
  MUX2_X2 U11102 ( .A(n7022), .B(n7021), .S(net366977), .Z(n7026) );
  NAND2_X2 U11103 ( .A1(daddr[30]), .A2(net368221), .ZN(n7031) );
  MUX2_X2 U11104 ( .A(regBoiz_regfile_0__2_), .B(regBoiz_regfile_1__2_), .S(
        net375713), .Z(n7033) );
  MUX2_X2 U11105 ( .A(regBoiz_regfile_2__2_), .B(regBoiz_regfile_3__2_), .S(
        net367025), .Z(n7032) );
  MUX2_X2 U11106 ( .A(n7033), .B(n7032), .S(net366977), .Z(n7037) );
  MUX2_X2 U11107 ( .A(regBoiz_regfile_4__2_), .B(regBoiz_regfile_5__2_), .S(
        net367027), .Z(n7035) );
  MUX2_X2 U11108 ( .A(regBoiz_regfile_6__2_), .B(regBoiz_regfile_7__2_), .S(
        net375717), .Z(n7034) );
  MUX2_X2 U11109 ( .A(n7035), .B(n7034), .S(net366977), .Z(n7036) );
  MUX2_X2 U11110 ( .A(n7037), .B(n7036), .S(net366933), .Z(n7045) );
  MUX2_X2 U11111 ( .A(regBoiz_regfile_8__2_), .B(regBoiz_regfile_9__2_), .S(
        net375713), .Z(n7039) );
  MUX2_X2 U11112 ( .A(regBoiz_regfile_10__2_), .B(regBoiz_regfile_11__2_), .S(
        net367029), .Z(n7038) );
  MUX2_X2 U11113 ( .A(n7039), .B(n7038), .S(net366977), .Z(n7043) );
  MUX2_X2 U11114 ( .A(regBoiz_regfile_12__2_), .B(regBoiz_regfile_13__2_), .S(
        net367023), .Z(n7041) );
  MUX2_X2 U11115 ( .A(regBoiz_regfile_14__2_), .B(regBoiz_regfile_15__2_), .S(
        net368800), .Z(n7040) );
  MUX2_X2 U11116 ( .A(n7041), .B(n7040), .S(net366977), .Z(n7042) );
  MUX2_X2 U11117 ( .A(n7043), .B(n7042), .S(net366933), .Z(n7044) );
  MUX2_X2 U11118 ( .A(n7045), .B(n7044), .S(net376330), .Z(n7061) );
  MUX2_X2 U11119 ( .A(regBoiz_regfile_16__2_), .B(regBoiz_regfile_17__2_), .S(
        net367029), .Z(n7047) );
  MUX2_X2 U11120 ( .A(regBoiz_regfile_18__2_), .B(regBoiz_regfile_19__2_), .S(
        net367027), .Z(n7046) );
  MUX2_X2 U11121 ( .A(n7047), .B(n7046), .S(net366987), .Z(n7051) );
  MUX2_X2 U11122 ( .A(regBoiz_regfile_20__2_), .B(regBoiz_regfile_21__2_), .S(
        net367031), .Z(n7049) );
  MUX2_X2 U11123 ( .A(regBoiz_regfile_22__2_), .B(regBoiz_regfile_23__2_), .S(
        net376223), .Z(n7048) );
  MUX2_X2 U11124 ( .A(n7049), .B(n7048), .S(net366977), .Z(n7050) );
  MUX2_X2 U11125 ( .A(n7051), .B(n7050), .S(net366939), .Z(n7059) );
  MUX2_X2 U11126 ( .A(regBoiz_regfile_24__2_), .B(regBoiz_regfile_25__2_), .S(
        net367025), .Z(n7053) );
  MUX2_X2 U11127 ( .A(regBoiz_regfile_26__2_), .B(regBoiz_regfile_27__2_), .S(
        net367019), .Z(n7052) );
  MUX2_X2 U11128 ( .A(n7053), .B(n7052), .S(net366977), .Z(n7057) );
  MUX2_X2 U11129 ( .A(regBoiz_regfile_28__2_), .B(regBoiz_regfile_29__2_), .S(
        net376222), .Z(n7055) );
  MUX2_X2 U11130 ( .A(regBoiz_regfile_30__2_), .B(n6311), .S(net375650), .Z(
        n7054) );
  MUX2_X2 U11131 ( .A(n7057), .B(n7056), .S(net366933), .Z(n7058) );
  MUX2_X2 U11132 ( .A(n7059), .B(n7058), .S(net376331), .Z(n7060) );
  NAND2_X2 U11133 ( .A1(daddr[29]), .A2(net368221), .ZN(n7062) );
  MUX2_X2 U11134 ( .A(regBoiz_regfile_0__3_), .B(regBoiz_regfile_1__3_), .S(
        net367031), .Z(n7064) );
  MUX2_X2 U11135 ( .A(regBoiz_regfile_2__3_), .B(regBoiz_regfile_3__3_), .S(
        net375718), .Z(n7063) );
  MUX2_X2 U11136 ( .A(n7064), .B(n7063), .S(net366977), .Z(n7068) );
  MUX2_X2 U11137 ( .A(regBoiz_regfile_4__3_), .B(regBoiz_regfile_5__3_), .S(
        net367027), .Z(n7066) );
  MUX2_X2 U11138 ( .A(regBoiz_regfile_6__3_), .B(regBoiz_regfile_7__3_), .S(
        net367029), .Z(n7065) );
  MUX2_X2 U11139 ( .A(n7066), .B(n7065), .S(net366977), .Z(n7067) );
  MUX2_X2 U11140 ( .A(n7068), .B(n7067), .S(net366933), .Z(n7076) );
  MUX2_X2 U11141 ( .A(regBoiz_regfile_8__3_), .B(regBoiz_regfile_9__3_), .S(
        net367029), .Z(n7070) );
  MUX2_X2 U11142 ( .A(regBoiz_regfile_10__3_), .B(regBoiz_regfile_11__3_), .S(
        net375717), .Z(n7069) );
  MUX2_X2 U11143 ( .A(n7070), .B(n7069), .S(net366977), .Z(n7074) );
  MUX2_X2 U11144 ( .A(regBoiz_regfile_12__3_), .B(regBoiz_regfile_13__3_), .S(
        net375718), .Z(n7072) );
  MUX2_X2 U11145 ( .A(n7072), .B(n7071), .S(net366977), .Z(n7073) );
  MUX2_X2 U11146 ( .A(n7074), .B(n7073), .S(net366919), .Z(n7075) );
  MUX2_X2 U11147 ( .A(n7076), .B(n7075), .S(net376331), .Z(n7092) );
  MUX2_X2 U11148 ( .A(regBoiz_regfile_16__3_), .B(regBoiz_regfile_24__3_), .S(
        net366899), .Z(n7078) );
  MUX2_X2 U11149 ( .A(regBoiz_regfile_18__3_), .B(regBoiz_regfile_26__3_), .S(
        net368781), .Z(n7077) );
  MUX2_X2 U11150 ( .A(n7078), .B(n7077), .S(net366979), .Z(n7082) );
  MUX2_X2 U11151 ( .A(regBoiz_regfile_20__3_), .B(regBoiz_regfile_28__3_), .S(
        net377166), .Z(n7080) );
  MUX2_X2 U11152 ( .A(regBoiz_regfile_22__3_), .B(n6464), .S(net376374), .Z(
        n7079) );
  MUX2_X2 U11153 ( .A(n7080), .B(n7079), .S(net366979), .Z(n7081) );
  MUX2_X2 U11154 ( .A(n7082), .B(n7081), .S(net378321), .Z(n7090) );
  MUX2_X2 U11155 ( .A(regBoiz_regfile_17__3_), .B(regBoiz_regfile_25__3_), .S(
        net366899), .Z(n7084) );
  MUX2_X2 U11156 ( .A(regBoiz_regfile_19__3_), .B(n6461), .S(net368781), .Z(
        n7083) );
  MUX2_X2 U11157 ( .A(n7084), .B(n7083), .S(net366979), .Z(n7088) );
  MUX2_X2 U11158 ( .A(n7086), .B(n7085), .S(net366979), .Z(n7087) );
  MUX2_X2 U11159 ( .A(n7088), .B(n7087), .S(net378321), .Z(n7089) );
  MUX2_X2 U11160 ( .A(n7090), .B(n7089), .S(net375718), .Z(n7091) );
  NAND2_X2 U11161 ( .A1(daddr[28]), .A2(net368221), .ZN(n9804) );
  MUX2_X2 U11162 ( .A(n7095), .B(n7094), .S(net366979), .Z(n7099) );
  MUX2_X2 U11163 ( .A(n7099), .B(n7098), .S(net366919), .Z(n7106) );
  MUX2_X2 U11164 ( .A(regBoiz_regfile_1__4_), .B(n6315), .S(net377464), .Z(
        n7100) );
  MUX2_X2 U11165 ( .A(n6313), .B(n6337), .S(n4978), .Z(n7102) );
  MUX2_X2 U11166 ( .A(regBoiz_regfile_16__4_), .B(regBoiz_regfile_24__4_), .S(
        net377166), .Z(n7108) );
  MUX2_X2 U11167 ( .A(n7112), .B(n7111), .S(net366939), .Z(n7118) );
  MUX2_X2 U11168 ( .A(n7114), .B(n7113), .S(net375527), .Z(n7116) );
  MUX2_X2 U11169 ( .A(n7120), .B(n7119), .S(n6784), .Z(n7121) );
  NAND2_X2 U11170 ( .A1(daddr[27]), .A2(net368221), .ZN(n9803) );
  MUX2_X2 U11171 ( .A(regBoiz_regfile_0__5_), .B(regBoiz_regfile_8__5_), .S(
        net368781), .Z(n7123) );
  MUX2_X2 U11172 ( .A(regBoiz_regfile_2__5_), .B(regBoiz_regfile_10__5_), .S(
        net377464), .Z(n7122) );
  MUX2_X2 U11173 ( .A(n7123), .B(n7122), .S(net366985), .Z(n7127) );
  MUX2_X2 U11174 ( .A(regBoiz_regfile_4__5_), .B(regBoiz_regfile_12__5_), .S(
        net369204), .Z(n7125) );
  MUX2_X2 U11175 ( .A(regBoiz_regfile_6__5_), .B(regBoiz_regfile_14__5_), .S(
        net376374), .Z(n7124) );
  MUX2_X2 U11176 ( .A(n7125), .B(n7124), .S(net366967), .Z(n7126) );
  MUX2_X2 U11177 ( .A(n7127), .B(n7126), .S(net366919), .Z(n7135) );
  MUX2_X2 U11178 ( .A(regBoiz_regfile_16__5_), .B(regBoiz_regfile_24__5_), .S(
        net377166), .Z(n7129) );
  MUX2_X2 U11179 ( .A(regBoiz_regfile_18__5_), .B(regBoiz_regfile_26__5_), .S(
        net366899), .Z(n7128) );
  MUX2_X2 U11180 ( .A(n7129), .B(n7128), .S(net366985), .Z(n7133) );
  MUX2_X2 U11181 ( .A(n7135), .B(n7134), .S(n6786), .Z(n7151) );
  MUX2_X2 U11182 ( .A(regBoiz_regfile_1__5_), .B(regBoiz_regfile_9__5_), .S(
        net369204), .Z(n7137) );
  MUX2_X2 U11183 ( .A(regBoiz_regfile_3__5_), .B(regBoiz_regfile_11__5_), .S(
        net377464), .Z(n7136) );
  MUX2_X2 U11184 ( .A(n7137), .B(n7136), .S(net366967), .Z(n7141) );
  MUX2_X2 U11185 ( .A(regBoiz_regfile_5__5_), .B(regBoiz_regfile_13__5_), .S(
        net377464), .Z(n7139) );
  MUX2_X2 U11186 ( .A(regBoiz_regfile_7__5_), .B(regBoiz_regfile_15__5_), .S(
        net377166), .Z(n7138) );
  MUX2_X2 U11187 ( .A(n7139), .B(n7138), .S(net366967), .Z(n7140) );
  MUX2_X2 U11188 ( .A(n7141), .B(n7140), .S(net378321), .Z(n7149) );
  MUX2_X2 U11189 ( .A(regBoiz_regfile_17__5_), .B(regBoiz_regfile_25__5_), .S(
        net366899), .Z(n7143) );
  MUX2_X2 U11190 ( .A(regBoiz_regfile_19__5_), .B(regBoiz_regfile_27__5_), .S(
        net369204), .Z(n7142) );
  MUX2_X2 U11191 ( .A(regBoiz_regfile_21__5_), .B(n6044), .S(net368770), .Z(
        n7145) );
  MUX2_X2 U11192 ( .A(regBoiz_regfile_23__5_), .B(regBoiz_regfile_31__5_), .S(
        net377166), .Z(n7144) );
  MUX2_X2 U11193 ( .A(n7149), .B(n7148), .S(n6784), .Z(n7150) );
  NAND2_X2 U11194 ( .A1(daddr[26]), .A2(net368221), .ZN(n9805) );
  MUX2_X2 U11195 ( .A(regBoiz_regfile_0__6_), .B(regBoiz_regfile_1__6_), .S(
        net367025), .Z(n7154) );
  MUX2_X2 U11196 ( .A(regBoiz_regfile_2__6_), .B(regBoiz_regfile_3__6_), .S(
        net367027), .Z(n7153) );
  MUX2_X2 U11197 ( .A(n7154), .B(n7153), .S(net366967), .Z(n7158) );
  MUX2_X2 U11198 ( .A(regBoiz_regfile_4__6_), .B(regBoiz_regfile_5__6_), .S(
        net375717), .Z(n7156) );
  MUX2_X2 U11199 ( .A(regBoiz_regfile_6__6_), .B(regBoiz_regfile_7__6_), .S(
        net367023), .Z(n7155) );
  MUX2_X2 U11200 ( .A(n7158), .B(n7157), .S(net378321), .Z(n7166) );
  MUX2_X2 U11201 ( .A(regBoiz_regfile_8__6_), .B(regBoiz_regfile_9__6_), .S(
        net375718), .Z(n7160) );
  MUX2_X2 U11202 ( .A(regBoiz_regfile_10__6_), .B(regBoiz_regfile_11__6_), .S(
        net367029), .Z(n7159) );
  MUX2_X2 U11203 ( .A(n7160), .B(n7159), .S(net366977), .Z(n7164) );
  MUX2_X2 U11204 ( .A(regBoiz_regfile_12__6_), .B(regBoiz_regfile_13__6_), .S(
        net367019), .Z(n7162) );
  MUX2_X2 U11205 ( .A(n7166), .B(n7165), .S(net375727), .Z(n7182) );
  MUX2_X2 U11206 ( .A(regBoiz_regfile_16__6_), .B(regBoiz_regfile_17__6_), .S(
        net367029), .Z(n7168) );
  MUX2_X2 U11207 ( .A(regBoiz_regfile_18__6_), .B(regBoiz_regfile_19__6_), .S(
        net367029), .Z(n7167) );
  MUX2_X2 U11208 ( .A(n7168), .B(n7167), .S(net375527), .Z(n7172) );
  MUX2_X2 U11209 ( .A(regBoiz_regfile_20__6_), .B(regBoiz_regfile_21__6_), .S(
        net367029), .Z(n7170) );
  MUX2_X2 U11210 ( .A(regBoiz_regfile_22__6_), .B(regBoiz_regfile_23__6_), .S(
        net375717), .Z(n7169) );
  MUX2_X2 U11211 ( .A(n7170), .B(n7169), .S(net366967), .Z(n7171) );
  MUX2_X2 U11212 ( .A(n7172), .B(n7171), .S(net366933), .Z(n7180) );
  MUX2_X2 U11213 ( .A(regBoiz_regfile_24__6_), .B(regBoiz_regfile_25__6_), .S(
        net367029), .Z(n7174) );
  MUX2_X2 U11214 ( .A(n7174), .B(n7173), .S(net366967), .Z(n7178) );
  MUX2_X2 U11215 ( .A(regBoiz_regfile_28__6_), .B(regBoiz_regfile_29__6_), .S(
        net367019), .Z(n7176) );
  MUX2_X2 U11216 ( .A(n7180), .B(n7179), .S(net375727), .Z(n7181) );
  NAND2_X2 U11217 ( .A1(daddr[25]), .A2(net368221), .ZN(n11769) );
  MUX2_X2 U11218 ( .A(regBoiz_regfile_0__7_), .B(regBoiz_regfile_1__7_), .S(
        net376222), .Z(n7185) );
  MUX2_X2 U11219 ( .A(regBoiz_regfile_2__7_), .B(regBoiz_regfile_3__7_), .S(
        net376223), .Z(n7184) );
  MUX2_X2 U11220 ( .A(n7185), .B(n7184), .S(net366967), .Z(n7189) );
  MUX2_X2 U11221 ( .A(regBoiz_regfile_4__7_), .B(regBoiz_regfile_5__7_), .S(
        net376222), .Z(n7187) );
  MUX2_X2 U11222 ( .A(regBoiz_regfile_6__7_), .B(n6307), .S(net367023), .Z(
        n7186) );
  MUX2_X2 U11223 ( .A(n7187), .B(n7186), .S(net366967), .Z(n7188) );
  MUX2_X2 U11224 ( .A(n7189), .B(n7188), .S(net366933), .Z(n7197) );
  MUX2_X2 U11225 ( .A(regBoiz_regfile_8__7_), .B(regBoiz_regfile_9__7_), .S(
        net367023), .Z(n7191) );
  MUX2_X2 U11226 ( .A(regBoiz_regfile_10__7_), .B(n6324), .S(net368800), .Z(
        n7190) );
  MUX2_X2 U11227 ( .A(n7191), .B(n7190), .S(net366967), .Z(n7195) );
  MUX2_X2 U11228 ( .A(regBoiz_regfile_12__7_), .B(n6309), .S(net376222), .Z(
        n7193) );
  MUX2_X2 U11229 ( .A(n7197), .B(n7196), .S(net375727), .Z(n7213) );
  MUX2_X2 U11230 ( .A(regBoiz_regfile_16__7_), .B(regBoiz_regfile_17__7_), .S(
        net376223), .Z(n7199) );
  MUX2_X2 U11231 ( .A(regBoiz_regfile_18__7_), .B(regBoiz_regfile_19__7_), .S(
        net376223), .Z(n7198) );
  MUX2_X2 U11232 ( .A(n7199), .B(n7198), .S(net366967), .Z(n7203) );
  MUX2_X2 U11233 ( .A(regBoiz_regfile_20__7_), .B(regBoiz_regfile_21__7_), .S(
        net367019), .Z(n7201) );
  MUX2_X2 U11234 ( .A(regBoiz_regfile_22__7_), .B(regBoiz_regfile_23__7_), .S(
        net367019), .Z(n7200) );
  MUX2_X2 U11235 ( .A(n7201), .B(n7200), .S(net366981), .Z(n7202) );
  MUX2_X2 U11236 ( .A(n7203), .B(n7202), .S(net378321), .Z(n7211) );
  MUX2_X2 U11237 ( .A(regBoiz_regfile_24__7_), .B(regBoiz_regfile_25__7_), .S(
        net376223), .Z(n7205) );
  MUX2_X2 U11238 ( .A(regBoiz_regfile_26__7_), .B(regBoiz_regfile_27__7_), .S(
        net367019), .Z(n7204) );
  MUX2_X2 U11239 ( .A(n7205), .B(n7204), .S(net366981), .Z(n7209) );
  MUX2_X2 U11240 ( .A(regBoiz_regfile_28__7_), .B(regBoiz_regfile_29__7_), .S(
        net376223), .Z(n7207) );
  MUX2_X2 U11241 ( .A(regBoiz_regfile_30__7_), .B(regBoiz_regfile_31__7_), .S(
        net367023), .Z(n7206) );
  MUX2_X2 U11242 ( .A(n7207), .B(n7206), .S(net366981), .Z(n7208) );
  MUX2_X2 U11243 ( .A(n7209), .B(n7208), .S(net366933), .Z(n7210) );
  NAND2_X2 U11244 ( .A1(daddr[24]), .A2(net368221), .ZN(n11726) );
  MUX2_X2 U11245 ( .A(regBoiz_regfile_0__8_), .B(regBoiz_regfile_1__8_), .S(
        net367023), .Z(n7216) );
  MUX2_X2 U11246 ( .A(regBoiz_regfile_2__8_), .B(regBoiz_regfile_3__8_), .S(
        net367019), .Z(n7215) );
  MUX2_X2 U11247 ( .A(n7216), .B(n7215), .S(net366981), .Z(n7220) );
  MUX2_X2 U11248 ( .A(regBoiz_regfile_4__8_), .B(regBoiz_regfile_5__8_), .S(
        net376222), .Z(n7218) );
  MUX2_X2 U11249 ( .A(regBoiz_regfile_6__8_), .B(regBoiz_regfile_7__8_), .S(
        net367023), .Z(n7217) );
  MUX2_X2 U11250 ( .A(n7218), .B(n7217), .S(net366981), .Z(n7219) );
  MUX2_X2 U11251 ( .A(n7220), .B(n7219), .S(net378321), .Z(n7228) );
  MUX2_X2 U11252 ( .A(regBoiz_regfile_8__8_), .B(regBoiz_regfile_9__8_), .S(
        net367023), .Z(n7222) );
  MUX2_X2 U11253 ( .A(regBoiz_regfile_10__8_), .B(regBoiz_regfile_11__8_), .S(
        net376223), .Z(n7221) );
  MUX2_X2 U11254 ( .A(n7222), .B(n7221), .S(net366981), .Z(n7226) );
  MUX2_X2 U11255 ( .A(regBoiz_regfile_12__8_), .B(regBoiz_regfile_13__8_), .S(
        net376223), .Z(n7224) );
  MUX2_X2 U11256 ( .A(n7228), .B(n7227), .S(n5242), .Z(n7229) );
  NAND2_X2 U11257 ( .A1(daddr[23]), .A2(net368221), .ZN(n9800) );
  MUX2_X2 U11258 ( .A(regBoiz_regfile_16__8_), .B(regBoiz_regfile_17__8_), .S(
        net376223), .Z(n7232) );
  MUX2_X2 U11259 ( .A(regBoiz_regfile_18__8_), .B(regBoiz_regfile_19__8_), .S(
        net367023), .Z(n7231) );
  MUX2_X2 U11260 ( .A(n7232), .B(n7231), .S(net366981), .Z(n7236) );
  MUX2_X2 U11261 ( .A(regBoiz_regfile_20__8_), .B(regBoiz_regfile_21__8_), .S(
        net376222), .Z(n7234) );
  MUX2_X2 U11262 ( .A(n7234), .B(n7233), .S(net366981), .Z(n7235) );
  MUX2_X2 U11263 ( .A(n7236), .B(n7235), .S(net366919), .Z(n7244) );
  MUX2_X2 U11264 ( .A(regBoiz_regfile_24__8_), .B(regBoiz_regfile_25__8_), .S(
        net367019), .Z(n7238) );
  MUX2_X2 U11265 ( .A(regBoiz_regfile_26__8_), .B(regBoiz_regfile_27__8_), .S(
        net367019), .Z(n7237) );
  MUX2_X2 U11266 ( .A(n7238), .B(n7237), .S(net366981), .Z(n7242) );
  MUX2_X2 U11267 ( .A(regBoiz_regfile_28__8_), .B(regBoiz_regfile_29__8_), .S(
        net376222), .Z(n7240) );
  MUX2_X2 U11268 ( .A(regBoiz_regfile_30__8_), .B(n6322), .S(net376223), .Z(
        n7239) );
  MUX2_X2 U11269 ( .A(n7244), .B(n7243), .S(net369204), .Z(n7245) );
  MUX2_X2 U11270 ( .A(regBoiz_regfile_0__9_), .B(regBoiz_regfile_8__9_), .S(
        net376077), .Z(n7248) );
  MUX2_X2 U11271 ( .A(regBoiz_regfile_2__9_), .B(regBoiz_regfile_10__9_), .S(
        net376331), .Z(n7247) );
  MUX2_X2 U11272 ( .A(n7248), .B(n7247), .S(net366981), .Z(n7252) );
  MUX2_X2 U11273 ( .A(regBoiz_regfile_4__9_), .B(regBoiz_regfile_12__9_), .S(
        net377464), .Z(n7250) );
  MUX2_X2 U11274 ( .A(regBoiz_regfile_6__9_), .B(n6445), .S(net376063), .Z(
        n7249) );
  MUX2_X2 U11275 ( .A(n7250), .B(n7249), .S(net366981), .Z(n7251) );
  MUX2_X2 U11276 ( .A(n7252), .B(n7251), .S(net366937), .Z(n7260) );
  MUX2_X2 U11277 ( .A(regBoiz_regfile_3__9_), .B(regBoiz_regfile_11__9_), .S(
        net368782), .Z(n7253) );
  MUX2_X2 U11278 ( .A(regBoiz_regfile_5__9_), .B(regBoiz_regfile_13__9_), .S(
        net368781), .Z(n7256) );
  MUX2_X2 U11279 ( .A(regBoiz_regfile_7__9_), .B(n6466), .S(net377464), .Z(
        n7255) );
  MUX2_X2 U11280 ( .A(regBoiz_regfile_16__9_), .B(regBoiz_regfile_24__9_), .S(
        net376330), .Z(n7262) );
  MUX2_X2 U11281 ( .A(regBoiz_regfile_18__9_), .B(n6449), .S(net377464), .Z(
        n7261) );
  MUX2_X2 U11282 ( .A(n7262), .B(n7261), .S(net366981), .Z(n7266) );
  MUX2_X2 U11283 ( .A(regBoiz_regfile_17__9_), .B(n6234), .S(net377464), .Z(
        n7268) );
  MUX2_X2 U11284 ( .A(n7268), .B(n7267), .S(net366981), .Z(n7272) );
  MUX2_X2 U11285 ( .A(regBoiz_regfile_21__9_), .B(n6468), .S(net377166), .Z(
        n7270) );
  NAND2_X2 U11286 ( .A1(daddr[22]), .A2(net368221), .ZN(n11719) );
  MUX2_X2 U11287 ( .A(regBoiz_regfile_0__10_), .B(regBoiz_regfile_8__10_), .S(
        net376063), .Z(n7279) );
  MUX2_X2 U11288 ( .A(regBoiz_regfile_2__10_), .B(regBoiz_regfile_10__10_), 
        .S(n5245), .Z(n7278) );
  MUX2_X2 U11289 ( .A(n7279), .B(n7278), .S(net366981), .Z(n7283) );
  MUX2_X2 U11290 ( .A(regBoiz_regfile_4__10_), .B(regBoiz_regfile_12__10_), 
        .S(net368782), .Z(n7281) );
  MUX2_X2 U11291 ( .A(regBoiz_regfile_6__10_), .B(n6396), .S(net368782), .Z(
        n7280) );
  MUX2_X2 U11292 ( .A(regBoiz_regfile_1__10_), .B(regBoiz_regfile_9__10_), .S(
        net375510), .Z(n7285) );
  MUX2_X2 U11293 ( .A(n7285), .B(n7284), .S(net366981), .Z(n7289) );
  MUX2_X2 U11294 ( .A(regBoiz_regfile_5__10_), .B(regBoiz_regfile_13__10_), 
        .S(net377464), .Z(n7287) );
  MUX2_X2 U11295 ( .A(regBoiz_regfile_7__10_), .B(n6447), .S(net366887), .Z(
        n7286) );
  MUX2_X2 U11296 ( .A(n7291), .B(n7290), .S(net376223), .Z(n7307) );
  MUX2_X2 U11297 ( .A(regBoiz_regfile_16__10_), .B(regBoiz_regfile_17__10_), 
        .S(net367019), .Z(n7293) );
  MUX2_X2 U11298 ( .A(regBoiz_regfile_18__10_), .B(regBoiz_regfile_19__10_), 
        .S(net376222), .Z(n7292) );
  MUX2_X2 U11299 ( .A(n7293), .B(n7292), .S(net366979), .Z(n7297) );
  MUX2_X2 U11300 ( .A(regBoiz_regfile_20__10_), .B(n6330), .S(net367023), .Z(
        n7295) );
  MUX2_X2 U11301 ( .A(regBoiz_regfile_22__10_), .B(n6451), .S(net367023), .Z(
        n7294) );
  MUX2_X2 U11302 ( .A(n7297), .B(n7296), .S(net366933), .Z(n7305) );
  MUX2_X2 U11303 ( .A(regBoiz_regfile_24__10_), .B(regBoiz_regfile_25__10_), 
        .S(net367019), .Z(n7299) );
  MUX2_X2 U11304 ( .A(regBoiz_regfile_26__10_), .B(n6453), .S(net376222), .Z(
        n7298) );
  MUX2_X2 U11305 ( .A(n7299), .B(n7298), .S(net366979), .Z(n7303) );
  MUX2_X2 U11306 ( .A(regBoiz_regfile_28__10_), .B(n6456), .S(net367019), .Z(
        n7301) );
  NAND2_X2 U11307 ( .A1(daddr[21]), .A2(net368221), .ZN(n11519) );
  NAND2_X2 U11308 ( .A1(n6787), .A2(net376330), .ZN(n7316) );
  INV_X4 U11309 ( .A(n7316), .ZN(n7312) );
  MUX2_X2 U11310 ( .A(regBoiz_regfile_24__11_), .B(regBoiz_regfile_25__11_), 
        .S(net367019), .Z(n7310) );
  MUX2_X2 U11311 ( .A(n7310), .B(n7309), .S(net366979), .Z(n7311) );
  NAND3_X2 U11312 ( .A1(n7312), .A2(n7311), .A3(net366953), .ZN(n7323) );
  MUX2_X2 U11313 ( .A(regBoiz_regfile_20__11_), .B(regBoiz_regfile_21__11_), 
        .S(net376223), .Z(n7314) );
  MUX2_X2 U11314 ( .A(regBoiz_regfile_22__11_), .B(regBoiz_regfile_23__11_), 
        .S(net376223), .Z(n7313) );
  MUX2_X2 U11315 ( .A(n7314), .B(n7313), .S(net366979), .Z(n7315) );
  MUX2_X2 U11316 ( .A(regBoiz_regfile_28__11_), .B(regBoiz_regfile_29__11_), 
        .S(net367019), .Z(n7318) );
  MUX2_X2 U11317 ( .A(regBoiz_regfile_30__11_), .B(regBoiz_regfile_31__11_), 
        .S(net367023), .Z(n7317) );
  MUX2_X2 U11318 ( .A(n7318), .B(n7317), .S(net366979), .Z(n7319) );
  MUX2_X2 U11319 ( .A(regBoiz_regfile_12__11_), .B(regBoiz_regfile_13__11_), 
        .S(net376223), .Z(n7325) );
  MUX2_X2 U11320 ( .A(regBoiz_regfile_14__11_), .B(regBoiz_regfile_15__11_), 
        .S(net376223), .Z(n7324) );
  MUX2_X2 U11321 ( .A(n7325), .B(n7324), .S(net366979), .Z(n7326) );
  NAND3_X2 U11322 ( .A1(net378321), .A2(n7326), .A3(n6794), .ZN(n7335) );
  MUX2_X2 U11323 ( .A(regBoiz_regfile_16__11_), .B(regBoiz_regfile_17__11_), 
        .S(net376222), .Z(n7328) );
  MUX2_X2 U11324 ( .A(n7328), .B(n7327), .S(net366979), .Z(n7329) );
  MUX2_X2 U11325 ( .A(regBoiz_regfile_8__11_), .B(regBoiz_regfile_9__11_), .S(
        net367023), .Z(n7331) );
  MUX2_X2 U11326 ( .A(n7331), .B(n7330), .S(net366977), .Z(n7332) );
  NAND3_X2 U11327 ( .A1(n7335), .A2(n7334), .A3(n7333), .ZN(n7347) );
  INV_X4 U11328 ( .A(n7336), .ZN(n7343) );
  MUX2_X2 U11329 ( .A(regBoiz_regfile_0__11_), .B(regBoiz_regfile_1__11_), .S(
        net376223), .Z(n7338) );
  MUX2_X2 U11330 ( .A(regBoiz_regfile_2__11_), .B(regBoiz_regfile_3__11_), .S(
        net376222), .Z(n7337) );
  MUX2_X2 U11331 ( .A(n7338), .B(n7337), .S(net366979), .Z(n7339) );
  MUX2_X2 U11332 ( .A(regBoiz_regfile_4__11_), .B(regBoiz_regfile_5__11_), .S(
        net367023), .Z(n7341) );
  MUX2_X2 U11333 ( .A(regBoiz_regfile_6__11_), .B(regBoiz_regfile_7__11_), .S(
        net376223), .Z(n7340) );
  MUX2_X2 U11334 ( .A(n7341), .B(n7340), .S(net366979), .Z(n7342) );
  NAND2_X2 U11335 ( .A1(daddr[20]), .A2(net368221), .ZN(n9815) );
  OAI22_X2 U11336 ( .A1(n7350), .A2(net375717), .B1(n7349), .B2(net367043), 
        .ZN(n7354) );
  MUX2_X2 U11337 ( .A(n7354), .B(n7353), .S(net366927), .Z(n7362) );
  MUX2_X2 U11338 ( .A(n7362), .B(n7361), .S(net368781), .Z(n7378) );
  AOI22_X2 U11339 ( .A1(regBoiz_regfile_20__12_), .A2(net367003), .B1(
        regBoiz_regfile_22__12_), .B2(net366985), .ZN(n7366) );
  AOI22_X2 U11340 ( .A1(regBoiz_regfile_21__12_), .A2(net367003), .B1(
        regBoiz_regfile_23__12_), .B2(net366985), .ZN(n7365) );
  OAI22_X2 U11341 ( .A1(n7366), .A2(net367027), .B1(n7365), .B2(net367041), 
        .ZN(n7367) );
  MUX2_X2 U11342 ( .A(n7368), .B(n7367), .S(net366927), .Z(n7376) );
  AOI22_X2 U11343 ( .A1(regBoiz_regfile_24__12_), .A2(net367003), .B1(
        regBoiz_regfile_26__12_), .B2(net366985), .ZN(n7370) );
  AOI22_X2 U11344 ( .A1(regBoiz_regfile_25__12_), .A2(net367003), .B1(
        regBoiz_regfile_27__12_), .B2(net366985), .ZN(n7369) );
  OAI22_X2 U11345 ( .A1(n7370), .A2(net367025), .B1(n7369), .B2(net367041), 
        .ZN(n7374) );
  OAI22_X2 U11346 ( .A1(n7372), .A2(net375717), .B1(n7371), .B2(net367041), 
        .ZN(n7373) );
  NAND2_X2 U11347 ( .A1(daddr[19]), .A2(net368221), .ZN(n9814) );
  OAI22_X2 U11348 ( .A1(n7381), .A2(net367027), .B1(n7380), .B2(net367041), 
        .ZN(n7385) );
  AOI22_X2 U11349 ( .A1(regBoiz_regfile_5__13_), .A2(net367003), .B1(
        regBoiz_regfile_7__13_), .B2(net366987), .ZN(n7382) );
  MUX2_X2 U11350 ( .A(n7385), .B(n7384), .S(net366927), .Z(n7393) );
  AOI22_X2 U11351 ( .A1(regBoiz_regfile_8__13_), .A2(net367001), .B1(
        regBoiz_regfile_10__13_), .B2(net366987), .ZN(n7387) );
  AOI22_X2 U11352 ( .A1(regBoiz_regfile_9__13_), .A2(net367003), .B1(
        regBoiz_regfile_11__13_), .B2(net366987), .ZN(n7386) );
  OAI22_X2 U11353 ( .A1(n7387), .A2(net367025), .B1(n7386), .B2(net367041), 
        .ZN(n7391) );
  AOI22_X2 U11354 ( .A1(regBoiz_regfile_12__13_), .A2(net367003), .B1(
        regBoiz_regfile_14__13_), .B2(net366987), .ZN(n7389) );
  AOI22_X2 U11355 ( .A1(regBoiz_regfile_13__13_), .A2(net367001), .B1(
        regBoiz_regfile_15__13_), .B2(net366987), .ZN(n7388) );
  OAI22_X2 U11356 ( .A1(n7389), .A2(net375718), .B1(n7388), .B2(net367041), 
        .ZN(n7390) );
  MUX2_X2 U11357 ( .A(n7391), .B(n7390), .S(net366919), .Z(n7392) );
  MUX2_X2 U11358 ( .A(n7393), .B(n7392), .S(net378488), .Z(n7408) );
  AOI22_X2 U11359 ( .A1(regBoiz_regfile_16__13_), .A2(net367001), .B1(
        regBoiz_regfile_18__13_), .B2(net366987), .ZN(n7395) );
  AOI22_X2 U11360 ( .A1(regBoiz_regfile_17__13_), .A2(net367001), .B1(
        regBoiz_regfile_19__13_), .B2(net366987), .ZN(n7394) );
  OAI22_X2 U11361 ( .A1(n7395), .A2(net375713), .B1(n7394), .B2(net367041), 
        .ZN(n7399) );
  AOI22_X2 U11362 ( .A1(regBoiz_regfile_20__13_), .A2(net367001), .B1(
        regBoiz_regfile_22__13_), .B2(net366987), .ZN(n7397) );
  AOI22_X2 U11363 ( .A1(regBoiz_regfile_21__13_), .A2(net367001), .B1(
        regBoiz_regfile_23__13_), .B2(net366987), .ZN(n7396) );
  OAI22_X2 U11364 ( .A1(n7397), .A2(net375713), .B1(n7396), .B2(net367041), 
        .ZN(n7398) );
  MUX2_X2 U11365 ( .A(n7399), .B(n7398), .S(net366927), .Z(n7406) );
  AOI22_X2 U11366 ( .A1(regBoiz_regfile_24__13_), .A2(net367001), .B1(
        regBoiz_regfile_26__13_), .B2(net366985), .ZN(n7401) );
  AOI22_X2 U11367 ( .A1(regBoiz_regfile_25__13_), .A2(net367001), .B1(
        regBoiz_regfile_27__13_), .B2(net366987), .ZN(n7400) );
  OAI22_X2 U11368 ( .A1(n7401), .A2(net367029), .B1(n7400), .B2(net367041), 
        .ZN(n7404) );
  OAI22_X2 U11369 ( .A1(net365830), .A2(net375718), .B1(n7402), .B2(net367043), 
        .ZN(n7403) );
  NAND2_X2 U11370 ( .A1(daddr[18]), .A2(net368221), .ZN(n9845) );
  NAND2_X2 U11371 ( .A1(regBoiz_regfile_6__14_), .A2(net366933), .ZN(n7410) );
  INV_X4 U11372 ( .A(n7410), .ZN(n7414) );
  NAND2_X2 U11373 ( .A1(regBoiz_regfile_4__14_), .A2(net366939), .ZN(n7411) );
  OAI211_X2 U11374 ( .C1(net378321), .C2(n5404), .A(n7411), .B(net367005), 
        .ZN(n7412) );
  OAI211_X2 U11375 ( .C1(n7414), .C2(n7413), .A(n7412), .B(net367043), .ZN(
        n7420) );
  NAND2_X2 U11376 ( .A1(regBoiz_regfile_5__14_), .A2(net378321), .ZN(n7415) );
  OAI211_X2 U11377 ( .C1(net366933), .C2(n5410), .A(n7415), .B(net367005), 
        .ZN(n7418) );
  NAND2_X2 U11378 ( .A1(regBoiz_regfile_7__14_), .A2(net366939), .ZN(n7416) );
  OAI211_X2 U11379 ( .C1(net366933), .C2(n5411), .A(net366987), .B(n7416), 
        .ZN(n7417) );
  NAND3_X2 U11380 ( .A1(net375713), .A2(n7418), .A3(n7417), .ZN(n7419) );
  NAND2_X2 U11381 ( .A1(n7420), .A2(n7419), .ZN(n7431) );
  NAND2_X2 U11382 ( .A1(regBoiz_regfile_12__14_), .A2(net366939), .ZN(n7421)
         );
  OAI211_X2 U11383 ( .C1(net366919), .C2(n5405), .A(n7421), .B(net367005), 
        .ZN(n7422) );
  OAI211_X2 U11384 ( .C1(n5447), .C2(n7423), .A(n7422), .B(net367043), .ZN(
        n7429) );
  NAND2_X2 U11385 ( .A1(regBoiz_regfile_13__14_), .A2(net366939), .ZN(n7424)
         );
  OAI211_X2 U11386 ( .C1(net366919), .C2(n5412), .A(n7424), .B(net367005), 
        .ZN(n7427) );
  NAND2_X2 U11387 ( .A1(regBoiz_regfile_15__14_), .A2(net366939), .ZN(n7425)
         );
  OAI211_X2 U11388 ( .C1(net366933), .C2(n5413), .A(net366987), .B(n7425), 
        .ZN(n7426) );
  NAND3_X2 U11389 ( .A1(net375650), .A2(n7427), .A3(n7426), .ZN(n7428) );
  NAND2_X2 U11390 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  MUX2_X2 U11391 ( .A(n7431), .B(n7430), .S(net378488), .Z(n7455) );
  NAND2_X2 U11392 ( .A1(regBoiz_regfile_22__14_), .A2(regBoiz_N12), .ZN(n7432)
         );
  INV_X4 U11393 ( .A(n7432), .ZN(n7436) );
  NAND2_X2 U11394 ( .A1(regBoiz_regfile_20__14_), .A2(net366937), .ZN(n7433)
         );
  OAI211_X2 U11395 ( .C1(net366933), .C2(n5406), .A(n7433), .B(net367005), 
        .ZN(n7434) );
  OAI211_X2 U11396 ( .C1(n7436), .C2(n7435), .A(n7434), .B(net367043), .ZN(
        n7442) );
  NAND2_X2 U11397 ( .A1(regBoiz_regfile_21__14_), .A2(net366937), .ZN(n7437)
         );
  OAI211_X2 U11398 ( .C1(net378321), .C2(n5414), .A(n7437), .B(net367005), 
        .ZN(n7440) );
  NAND2_X2 U11399 ( .A1(regBoiz_regfile_23__14_), .A2(net366937), .ZN(n7438)
         );
  OAI211_X2 U11400 ( .C1(net366933), .C2(n5415), .A(net366987), .B(n7438), 
        .ZN(n7439) );
  NAND3_X2 U11401 ( .A1(net367031), .A2(n7440), .A3(n7439), .ZN(n7441) );
  NAND2_X2 U11402 ( .A1(n7442), .A2(n7441), .ZN(n7453) );
  OAI211_X2 U11403 ( .C1(net366933), .C2(n5407), .A(n7443), .B(net367005), 
        .ZN(n7444) );
  OAI211_X2 U11404 ( .C1(n5448), .C2(n7445), .A(n7444), .B(net367043), .ZN(
        n7451) );
  NAND2_X2 U11405 ( .A1(regBoiz_regfile_29__14_), .A2(net366939), .ZN(n7446)
         );
  OAI211_X2 U11406 ( .C1(net366933), .C2(n5416), .A(n7446), .B(net367005), 
        .ZN(n7449) );
  OAI211_X2 U11407 ( .C1(net366933), .C2(n5417), .A(net366987), .B(n7447), 
        .ZN(n7448) );
  NAND3_X2 U11408 ( .A1(net375718), .A2(n7449), .A3(n7448), .ZN(n7450) );
  NAND2_X2 U11409 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  MUX2_X2 U11410 ( .A(n7455), .B(n7454), .S(n6785), .Z(n7456) );
  NAND2_X2 U11411 ( .A1(daddr[17]), .A2(net368221), .ZN(n9844) );
  INV_X4 U11412 ( .A(n9882), .ZN(n7483) );
  NAND3_X4 U11413 ( .A1(n7464), .A2(n7463), .A3(n7483), .ZN(n7475) );
  NAND2_X2 U11414 ( .A1(net369200), .A2(net375717), .ZN(n9880) );
  NAND3_X4 U11415 ( .A1(n7468), .A2(n7467), .A3(n7557), .ZN(n7474) );
  NAND4_X2 U11416 ( .A1(n7476), .A2(n7475), .A3(n7474), .A4(n7473), .ZN(n7499)
         );
  NOR2_X4 U11417 ( .A1(net366923), .A2(n5527), .ZN(n7477) );
  OAI21_X4 U11418 ( .B1(n5428), .B2(n7477), .A(net366999), .ZN(n7480) );
  NOR2_X4 U11419 ( .A1(net366923), .A2(n5528), .ZN(n7478) );
  OAI21_X4 U11420 ( .B1(n5429), .B2(n7478), .A(net366967), .ZN(n7479) );
  NAND3_X4 U11421 ( .A1(n7480), .A2(n7479), .A3(net365399), .ZN(n7497) );
  NOR2_X4 U11422 ( .A1(net366923), .A2(n5541), .ZN(n7481) );
  OAI21_X4 U11423 ( .B1(n5434), .B2(n7481), .A(net366999), .ZN(n7485) );
  NOR2_X4 U11424 ( .A1(net366923), .A2(n5542), .ZN(n7482) );
  OAI21_X4 U11425 ( .B1(n5435), .B2(n7482), .A(net366967), .ZN(n7484) );
  NAND3_X4 U11426 ( .A1(n7485), .A2(n7484), .A3(n7483), .ZN(n7496) );
  NOR2_X4 U11427 ( .A1(net366923), .A2(n5543), .ZN(n7486) );
  OAI21_X4 U11428 ( .B1(n5436), .B2(n7486), .A(net366999), .ZN(n7489) );
  NOR2_X4 U11429 ( .A1(net366925), .A2(n5544), .ZN(n7487) );
  NAND3_X4 U11430 ( .A1(n7489), .A2(n7488), .A3(n7557), .ZN(n7495) );
  NOR2_X4 U11431 ( .A1(net366923), .A2(n5529), .ZN(n7490) );
  OAI21_X4 U11432 ( .B1(n5430), .B2(n7490), .A(net366999), .ZN(n7493) );
  NOR2_X4 U11433 ( .A1(net366921), .A2(n5530), .ZN(n7491) );
  NAND3_X4 U11434 ( .A1(n7493), .A2(n7492), .A3(n6054), .ZN(n7494) );
  NAND4_X2 U11435 ( .A1(n7497), .A2(n7496), .A3(n7495), .A4(n7494), .ZN(n7498)
         );
  MUX2_X2 U11436 ( .A(n7499), .B(n7498), .S(n6784), .Z(n7501) );
  NAND2_X2 U11437 ( .A1(daddr[16]), .A2(net368221), .ZN(n7500) );
  MUX2_X2 U11438 ( .A(regBoiz_regfile_0__16_), .B(regBoiz_regfile_8__16_), .S(
        net366899), .Z(n7503) );
  MUX2_X2 U11439 ( .A(n7503), .B(n7502), .S(net366969), .Z(n7507) );
  MUX2_X2 U11440 ( .A(regBoiz_regfile_4__16_), .B(regBoiz_regfile_12__16_), 
        .S(net369200), .Z(n7505) );
  MUX2_X2 U11441 ( .A(n7507), .B(n7506), .S(net366919), .Z(n11052) );
  NAND2_X2 U11442 ( .A1(n6531), .A2(n11052), .ZN(n7530) );
  MUX2_X2 U11443 ( .A(regBoiz_regfile_16__16_), .B(regBoiz_regfile_24__16_), 
        .S(net376063), .Z(n7509) );
  MUX2_X2 U11444 ( .A(n7509), .B(n7508), .S(net366969), .Z(n7513) );
  MUX2_X2 U11445 ( .A(regBoiz_regfile_20__16_), .B(regBoiz_regfile_28__16_), 
        .S(net366887), .Z(n7511) );
  MUX2_X2 U11446 ( .A(regBoiz_regfile_22__16_), .B(regBoiz_regfile_30__16_), 
        .S(net377109), .Z(n7510) );
  MUX2_X2 U11447 ( .A(regBoiz_regfile_17__16_), .B(regBoiz_regfile_25__16_), 
        .S(net368782), .Z(n7516) );
  MUX2_X2 U11448 ( .A(regBoiz_regfile_19__16_), .B(regBoiz_regfile_27__16_), 
        .S(net366887), .Z(n7515) );
  MUX2_X2 U11449 ( .A(n7516), .B(n7515), .S(net366969), .Z(n7520) );
  MUX2_X2 U11450 ( .A(regBoiz_regfile_21__16_), .B(regBoiz_regfile_29__16_), 
        .S(net376374), .Z(n7518) );
  MUX2_X2 U11451 ( .A(regBoiz_regfile_23__16_), .B(n6022), .S(net375510), .Z(
        n7517) );
  MUX2_X2 U11452 ( .A(n7518), .B(n7517), .S(net366969), .Z(n7519) );
  MUX2_X2 U11453 ( .A(n7520), .B(n7519), .S(net366919), .Z(n9819) );
  NAND2_X2 U11454 ( .A1(net375713), .A2(n6794), .ZN(n9823) );
  INV_X4 U11455 ( .A(n9823), .ZN(n11053) );
  MUX2_X2 U11456 ( .A(regBoiz_regfile_1__16_), .B(regBoiz_regfile_9__16_), .S(
        net377166), .Z(n7523) );
  MUX2_X2 U11457 ( .A(regBoiz_regfile_3__16_), .B(regBoiz_regfile_11__16_), 
        .S(net378494), .Z(n7522) );
  MUX2_X2 U11458 ( .A(n7523), .B(n7522), .S(net366969), .Z(n7527) );
  MUX2_X2 U11459 ( .A(regBoiz_regfile_5__16_), .B(regBoiz_regfile_13__16_), 
        .S(net368781), .Z(n7525) );
  MUX2_X2 U11460 ( .A(n7527), .B(n7526), .S(net366933), .Z(n11054) );
  NAND3_X2 U11461 ( .A1(n7530), .A2(n7529), .A3(n7528), .ZN(n7531) );
  NAND2_X2 U11462 ( .A1(daddr[15]), .A2(net368221), .ZN(n11180) );
  NAND2_X2 U11463 ( .A1(daddr[14]), .A2(net368221), .ZN(n9833) );
  MUX2_X2 U11464 ( .A(regBoiz_regfile_0__17_), .B(regBoiz_regfile_16__17_), 
        .S(n6786), .Z(n7533) );
  MUX2_X2 U11465 ( .A(regBoiz_regfile_2__17_), .B(regBoiz_regfile_18__17_), 
        .S(n5093), .Z(n7532) );
  MUX2_X2 U11466 ( .A(n7533), .B(n7532), .S(net366969), .Z(n7535) );
  NOR2_X4 U11467 ( .A1(net366921), .A2(net368782), .ZN(n8039) );
  NAND2_X2 U11468 ( .A1(n8039), .A2(net367043), .ZN(n7534) );
  NOR2_X4 U11469 ( .A1(n7535), .A2(n7534), .ZN(n7541) );
  MUX2_X2 U11470 ( .A(regBoiz_regfile_4__17_), .B(regBoiz_regfile_20__17_), 
        .S(n6785), .Z(n7537) );
  MUX2_X2 U11471 ( .A(regBoiz_regfile_6__17_), .B(regBoiz_regfile_22__17_), 
        .S(n6785), .Z(n7536) );
  MUX2_X2 U11472 ( .A(n7537), .B(n7536), .S(net366969), .Z(n7539) );
  NAND2_X2 U11473 ( .A1(n7670), .A2(net367043), .ZN(n7538) );
  NOR2_X4 U11474 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  NOR2_X4 U11475 ( .A1(n7541), .A2(n7540), .ZN(n9831) );
  MUX2_X2 U11476 ( .A(regBoiz_regfile_1__17_), .B(regBoiz_regfile_17__17_), 
        .S(n6786), .Z(n7543) );
  MUX2_X2 U11477 ( .A(regBoiz_regfile_3__17_), .B(regBoiz_regfile_19__17_), 
        .S(n6782), .Z(n7542) );
  MUX2_X2 U11478 ( .A(n7543), .B(n7542), .S(net366969), .Z(n7547) );
  NOR2_X4 U11479 ( .A1(net366921), .A2(net369316), .ZN(n8025) );
  MUX2_X2 U11480 ( .A(regBoiz_regfile_8__17_), .B(regBoiz_regfile_24__17_), 
        .S(n6784), .Z(n7545) );
  MUX2_X2 U11481 ( .A(regBoiz_regfile_10__17_), .B(regBoiz_regfile_26__17_), 
        .S(n6782), .Z(n7544) );
  MUX2_X2 U11482 ( .A(regBoiz_regfile_12__17_), .B(regBoiz_regfile_28__17_), 
        .S(n6784), .Z(n7549) );
  MUX2_X2 U11483 ( .A(regBoiz_regfile_14__17_), .B(regBoiz_regfile_30__17_), 
        .S(n6786), .Z(n7548) );
  MUX2_X2 U11484 ( .A(n7549), .B(n7548), .S(net366971), .Z(n7550) );
  NAND2_X2 U11485 ( .A1(n9855), .A2(n7550), .ZN(n7563) );
  MUX2_X2 U11486 ( .A(regBoiz_regfile_5__17_), .B(regBoiz_regfile_21__17_), 
        .S(n6784), .Z(n7552) );
  MUX2_X2 U11487 ( .A(regBoiz_regfile_7__17_), .B(regBoiz_regfile_23__17_), 
        .S(n6784), .Z(n7551) );
  MUX2_X2 U11488 ( .A(n7552), .B(n7551), .S(net366969), .Z(n7556) );
  MUX2_X2 U11489 ( .A(regBoiz_regfile_9__17_), .B(regBoiz_regfile_25__17_), 
        .S(n6786), .Z(n7554) );
  MUX2_X2 U11490 ( .A(regBoiz_regfile_11__17_), .B(regBoiz_regfile_27__17_), 
        .S(n6785), .Z(n7553) );
  MUX2_X2 U11491 ( .A(regBoiz_regfile_13__17_), .B(regBoiz_regfile_29__17_), 
        .S(n6785), .Z(n7559) );
  MUX2_X2 U11492 ( .A(regBoiz_regfile_15__17_), .B(regBoiz_regfile_31__17_), 
        .S(n6784), .Z(n7558) );
  MUX2_X2 U11493 ( .A(n7559), .B(n7558), .S(net366971), .Z(n7560) );
  NAND3_X4 U11494 ( .A1(n9832), .A2(net362297), .A3(n9831), .ZN(n7565) );
  MUX2_X2 U11495 ( .A(regBoiz_regfile_4__18_), .B(regBoiz_regfile_20__18_), 
        .S(n6786), .Z(n7567) );
  MUX2_X2 U11496 ( .A(regBoiz_regfile_6__18_), .B(regBoiz_regfile_22__18_), 
        .S(n5107), .Z(n7566) );
  MUX2_X2 U11497 ( .A(n7567), .B(n7566), .S(net366971), .Z(n7573) );
  MUX2_X2 U11498 ( .A(regBoiz_regfile_0__18_), .B(regBoiz_regfile_16__18_), 
        .S(n6785), .Z(n7569) );
  MUX2_X2 U11499 ( .A(regBoiz_regfile_2__18_), .B(regBoiz_regfile_18__18_), 
        .S(n6784), .Z(n7568) );
  MUX2_X2 U11500 ( .A(n7569), .B(n7568), .S(net366971), .Z(n7571) );
  NAND2_X2 U11501 ( .A1(n8039), .A2(net367043), .ZN(n7570) );
  MUX2_X2 U11502 ( .A(regBoiz_regfile_1__18_), .B(regBoiz_regfile_17__18_), 
        .S(n6785), .Z(n7576) );
  MUX2_X2 U11503 ( .A(regBoiz_regfile_3__18_), .B(regBoiz_regfile_19__18_), 
        .S(n6784), .Z(n7575) );
  MUX2_X2 U11504 ( .A(n7576), .B(n7575), .S(net366971), .Z(n7580) );
  MUX2_X2 U11505 ( .A(regBoiz_regfile_8__18_), .B(regBoiz_regfile_24__18_), 
        .S(n6786), .Z(n7578) );
  MUX2_X2 U11506 ( .A(regBoiz_regfile_10__18_), .B(regBoiz_regfile_26__18_), 
        .S(n6786), .Z(n7577) );
  MUX2_X2 U11507 ( .A(regBoiz_regfile_12__18_), .B(regBoiz_regfile_28__18_), 
        .S(n6786), .Z(n7582) );
  MUX2_X2 U11508 ( .A(regBoiz_regfile_14__18_), .B(regBoiz_regfile_30__18_), 
        .S(n6785), .Z(n7581) );
  MUX2_X2 U11509 ( .A(n7582), .B(n7581), .S(net366971), .Z(n7583) );
  NAND2_X2 U11510 ( .A1(n9855), .A2(n7583), .ZN(n7595) );
  MUX2_X2 U11511 ( .A(regBoiz_regfile_5__18_), .B(regBoiz_regfile_21__18_), 
        .S(n6786), .Z(n7585) );
  MUX2_X2 U11512 ( .A(regBoiz_regfile_7__18_), .B(regBoiz_regfile_23__18_), 
        .S(n6785), .Z(n7584) );
  MUX2_X2 U11513 ( .A(n7585), .B(n7584), .S(net366971), .Z(n7589) );
  MUX2_X2 U11514 ( .A(regBoiz_regfile_9__18_), .B(regBoiz_regfile_25__18_), 
        .S(n6785), .Z(n7587) );
  MUX2_X2 U11515 ( .A(n7587), .B(n7586), .S(net366971), .Z(n7588) );
  MUX2_X2 U11516 ( .A(regBoiz_regfile_13__18_), .B(regBoiz_regfile_29__18_), 
        .S(n6784), .Z(n7591) );
  MUX2_X2 U11517 ( .A(regBoiz_regfile_15__18_), .B(regBoiz_regfile_31__18_), 
        .S(n6786), .Z(n7590) );
  NAND3_X4 U11518 ( .A1(n9830), .A2(net362297), .A3(n9829), .ZN(n7597) );
  MUX2_X2 U11519 ( .A(regBoiz_regfile_13__19_), .B(regBoiz_regfile_29__19_), 
        .S(n6786), .Z(n7599) );
  MUX2_X2 U11520 ( .A(regBoiz_regfile_15__19_), .B(regBoiz_regfile_31__19_), 
        .S(n6784), .Z(n7598) );
  MUX2_X2 U11521 ( .A(regBoiz_regfile_1__19_), .B(regBoiz_regfile_17__19_), 
        .S(n6785), .Z(n7602) );
  MUX2_X2 U11522 ( .A(regBoiz_regfile_3__19_), .B(regBoiz_regfile_19__19_), 
        .S(n6784), .Z(n7601) );
  MUX2_X2 U11523 ( .A(n7602), .B(n7601), .S(net366971), .Z(n7603) );
  NAND2_X2 U11524 ( .A1(n8039), .A2(n7603), .ZN(n7612) );
  MUX2_X2 U11525 ( .A(regBoiz_regfile_5__19_), .B(regBoiz_regfile_21__19_), 
        .S(n6784), .Z(n7605) );
  MUX2_X2 U11526 ( .A(regBoiz_regfile_7__19_), .B(regBoiz_regfile_23__19_), 
        .S(n6784), .Z(n7604) );
  MUX2_X2 U11527 ( .A(n7605), .B(n7604), .S(net366971), .Z(n7606) );
  NAND2_X2 U11528 ( .A1(n7670), .A2(n7606), .ZN(n7611) );
  MUX2_X2 U11529 ( .A(regBoiz_regfile_9__19_), .B(regBoiz_regfile_25__19_), 
        .S(n6786), .Z(n7608) );
  MUX2_X2 U11530 ( .A(regBoiz_regfile_11__19_), .B(regBoiz_regfile_27__19_), 
        .S(n6785), .Z(n7607) );
  MUX2_X2 U11531 ( .A(n7608), .B(n7607), .S(net366971), .Z(n7609) );
  NAND2_X2 U11532 ( .A1(net365293), .A2(n7609), .ZN(n7610) );
  NAND4_X2 U11533 ( .A1(n7613), .A2(n7612), .A3(n7611), .A4(n7610), .ZN(n7638)
         );
  NAND2_X2 U11534 ( .A1(regBoiz_regfile_6__19_), .A2(net366933), .ZN(n7614) );
  NAND2_X2 U11535 ( .A1(regBoiz_regfile_22__19_), .A2(net366933), .ZN(n7616)
         );
  OAI211_X2 U11536 ( .C1(net366933), .C2(n5566), .A(n6787), .B(n7616), .ZN(
        n7622) );
  NAND2_X2 U11537 ( .A1(regBoiz_regfile_4__19_), .A2(net366933), .ZN(n7619) );
  AOI22_X2 U11538 ( .A1(n7623), .A2(n7622), .B1(n7621), .B2(n7620), .ZN(n7635)
         );
  NAND2_X2 U11539 ( .A1(regBoiz_regfile_14__19_), .A2(net366919), .ZN(n7624)
         );
  AOI21_X4 U11540 ( .B1(n7625), .B2(n7624), .A(net366999), .ZN(n7633) );
  NAND2_X2 U11541 ( .A1(regBoiz_regfile_30__19_), .A2(net366919), .ZN(n7626)
         );
  OAI211_X2 U11542 ( .C1(net366933), .C2(n5567), .A(n6787), .B(n7626), .ZN(
        n7632) );
  NAND2_X2 U11543 ( .A1(regBoiz_regfile_28__19_), .A2(net366919), .ZN(n7627)
         );
  NAND2_X2 U11544 ( .A1(regBoiz_regfile_12__19_), .A2(net366919), .ZN(n7629)
         );
  OAI211_X2 U11545 ( .C1(net366933), .C2(n5568), .A(n6794), .B(n7629), .ZN(
        n7630) );
  AOI22_X2 U11546 ( .A1(n7633), .A2(n7632), .B1(n7631), .B2(n7630), .ZN(n7634)
         );
  MUX2_X2 U11547 ( .A(n7635), .B(n7634), .S(net368781), .Z(n7636) );
  NAND2_X2 U11548 ( .A1(n7636), .A2(net367045), .ZN(n7637) );
  MUX2_X2 U11549 ( .A(regBoiz_regfile_9__20_), .B(regBoiz_regfile_25__20_), 
        .S(n6784), .Z(n7641) );
  MUX2_X2 U11550 ( .A(regBoiz_regfile_11__20_), .B(regBoiz_regfile_27__20_), 
        .S(n6786), .Z(n7640) );
  MUX2_X2 U11551 ( .A(n7641), .B(n7640), .S(net366971), .Z(n7642) );
  NAND3_X2 U11552 ( .A1(net375713), .A2(n7642), .A3(net365293), .ZN(n7651) );
  MUX2_X2 U11553 ( .A(regBoiz_regfile_5__20_), .B(regBoiz_regfile_21__20_), 
        .S(n6784), .Z(n7644) );
  MUX2_X2 U11554 ( .A(regBoiz_regfile_7__20_), .B(regBoiz_regfile_23__20_), 
        .S(n6785), .Z(n7643) );
  MUX2_X2 U11555 ( .A(n7644), .B(n7643), .S(net366971), .Z(n7645) );
  MUX2_X2 U11556 ( .A(regBoiz_regfile_13__20_), .B(regBoiz_regfile_29__20_), 
        .S(n6784), .Z(n7647) );
  MUX2_X2 U11557 ( .A(regBoiz_regfile_15__20_), .B(regBoiz_regfile_31__20_), 
        .S(n6785), .Z(n7646) );
  MUX2_X2 U11558 ( .A(regBoiz_regfile_8__20_), .B(regBoiz_regfile_24__20_), 
        .S(n6785), .Z(n7653) );
  MUX2_X2 U11559 ( .A(regBoiz_regfile_10__20_), .B(regBoiz_regfile_26__20_), 
        .S(n6784), .Z(n7652) );
  MUX2_X2 U11560 ( .A(n7653), .B(n7652), .S(net366971), .Z(n7654) );
  NAND2_X2 U11561 ( .A1(n8025), .A2(n7654), .ZN(n7663) );
  MUX2_X2 U11562 ( .A(regBoiz_regfile_1__20_), .B(regBoiz_regfile_17__20_), 
        .S(n6786), .Z(n7656) );
  MUX2_X2 U11563 ( .A(n7656), .B(n7655), .S(net366971), .Z(n7657) );
  NAND2_X2 U11564 ( .A1(n8039), .A2(n7657), .ZN(n7662) );
  MUX2_X2 U11565 ( .A(regBoiz_regfile_12__20_), .B(regBoiz_regfile_28__20_), 
        .S(n6785), .Z(n7659) );
  MUX2_X2 U11566 ( .A(n7659), .B(n7658), .S(net366971), .Z(n7660) );
  NAND2_X2 U11567 ( .A1(n9855), .A2(n7660), .ZN(n7661) );
  NAND3_X2 U11568 ( .A1(n7663), .A2(n7662), .A3(n7661), .ZN(n7676) );
  MUX2_X2 U11569 ( .A(regBoiz_regfile_0__20_), .B(regBoiz_regfile_16__20_), 
        .S(n6782), .Z(n7665) );
  MUX2_X2 U11570 ( .A(regBoiz_regfile_2__20_), .B(regBoiz_regfile_18__20_), 
        .S(n6789), .Z(n7664) );
  MUX2_X2 U11571 ( .A(n7665), .B(n7664), .S(net366973), .Z(n7667) );
  NAND2_X2 U11572 ( .A1(n8039), .A2(net367043), .ZN(n7666) );
  NOR2_X4 U11573 ( .A1(n7667), .A2(n7666), .ZN(n7674) );
  MUX2_X2 U11574 ( .A(regBoiz_regfile_4__20_), .B(regBoiz_regfile_20__20_), 
        .S(n6782), .Z(n7669) );
  MUX2_X2 U11575 ( .A(regBoiz_regfile_6__20_), .B(regBoiz_regfile_22__20_), 
        .S(n6370), .Z(n7668) );
  MUX2_X2 U11576 ( .A(n7669), .B(n7668), .S(net366973), .Z(n7672) );
  NAND2_X2 U11577 ( .A1(n7670), .A2(net367043), .ZN(n7671) );
  NOR2_X4 U11578 ( .A1(n7672), .A2(n7671), .ZN(n7673) );
  NOR3_X4 U11579 ( .A1(net368548), .A2(n7674), .A3(n7673), .ZN(n7675) );
  OAI21_X4 U11580 ( .B1(n7677), .B2(n7676), .A(n7675), .ZN(n9895) );
  NAND2_X2 U11581 ( .A1(daddr[11]), .A2(net368223), .ZN(n9894) );
  NOR2_X4 U11582 ( .A1(net366921), .A2(n5545), .ZN(n7679) );
  NAND2_X2 U11583 ( .A1(regBoiz_regfile_13__21_), .A2(net366933), .ZN(n7682)
         );
  INV_X4 U11584 ( .A(n7682), .ZN(n7684) );
  NOR2_X4 U11585 ( .A1(net366921), .A2(n5547), .ZN(n7685) );
  NAND2_X2 U11586 ( .A1(regBoiz_regfile_31__21_), .A2(net366919), .ZN(n7690)
         );
  INV_X4 U11587 ( .A(n7690), .ZN(n7692) );
  NOR2_X4 U11588 ( .A1(net366921), .A2(n5549), .ZN(n7691) );
  NAND3_X4 U11589 ( .A1(n7698), .A2(n7697), .A3(n7696), .ZN(n7736) );
  NOR2_X4 U11590 ( .A1(net366921), .A2(n5396), .ZN(n7700) );
  NAND2_X2 U11591 ( .A1(regBoiz_regfile_23__21_), .A2(net366919), .ZN(n7705)
         );
  INV_X4 U11592 ( .A(n7705), .ZN(n7707) );
  NOR2_X4 U11593 ( .A1(net366921), .A2(n5402), .ZN(n7706) );
  NAND2_X2 U11594 ( .A1(net366987), .A2(net375929), .ZN(n8134) );
  INV_X4 U11595 ( .A(n8134), .ZN(n8147) );
  NAND2_X2 U11596 ( .A1(regBoiz_regfile_14__21_), .A2(net366919), .ZN(n7710)
         );
  INV_X4 U11597 ( .A(n7710), .ZN(n7712) );
  NOR2_X4 U11598 ( .A1(net366921), .A2(n5532), .ZN(n7711) );
  NOR2_X4 U11599 ( .A1(net366921), .A2(n5397), .ZN(n7713) );
  INV_X4 U11600 ( .A(net365399), .ZN(net364906) );
  NAND4_X2 U11601 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(net364906), .ZN(
        n7735) );
  NAND2_X2 U11602 ( .A1(regBoiz_regfile_22__21_), .A2(net366919), .ZN(n7721)
         );
  INV_X4 U11603 ( .A(n7721), .ZN(n7723) );
  NOR2_X4 U11604 ( .A1(net366921), .A2(n5534), .ZN(n7722) );
  NAND2_X2 U11605 ( .A1(regBoiz_regfile_4__21_), .A2(net366919), .ZN(n7726) );
  INV_X4 U11606 ( .A(n7726), .ZN(n7728) );
  NOR2_X4 U11607 ( .A1(net366921), .A2(n5535), .ZN(n7727) );
  NOR2_X4 U11608 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  OAI21_X4 U11609 ( .B1(n7736), .B2(n7735), .A(n7734), .ZN(net363047) );
  NAND2_X2 U11610 ( .A1(daddr[10]), .A2(net362342), .ZN(net363049) );
  NOR2_X4 U11611 ( .A1(net366923), .A2(n6782), .ZN(n9846) );
  MUX2_X2 U11612 ( .A(regBoiz_regfile_0__22_), .B(regBoiz_regfile_8__22_), .S(
        net366899), .Z(n7738) );
  MUX2_X2 U11613 ( .A(regBoiz_regfile_2__22_), .B(regBoiz_regfile_10__22_), 
        .S(net377166), .Z(n7737) );
  MUX2_X2 U11614 ( .A(n7738), .B(n7737), .S(net366973), .Z(n7739) );
  INV_X4 U11615 ( .A(n7739), .ZN(n9869) );
  MUX2_X2 U11616 ( .A(regBoiz_regfile_4__22_), .B(regBoiz_regfile_12__22_), 
        .S(net376374), .Z(n7741) );
  MUX2_X2 U11617 ( .A(regBoiz_regfile_6__22_), .B(regBoiz_regfile_14__22_), 
        .S(net376374), .Z(n7740) );
  MUX2_X2 U11618 ( .A(n7741), .B(n7740), .S(net366973), .Z(n9866) );
  NAND2_X2 U11619 ( .A1(net366919), .A2(n6795), .ZN(n9848) );
  MUX2_X2 U11620 ( .A(regBoiz_regfile_5__22_), .B(regBoiz_regfile_13__22_), 
        .S(net369204), .Z(n7744) );
  MUX2_X2 U11621 ( .A(regBoiz_regfile_7__22_), .B(regBoiz_regfile_15__22_), 
        .S(n5245), .Z(n7743) );
  MUX2_X2 U11622 ( .A(regBoiz_regfile_22__22_), .B(regBoiz_regfile_30__22_), 
        .S(net376077), .Z(n7746) );
  NAND2_X2 U11623 ( .A1(net366987), .A2(n7746), .ZN(n9857) );
  MUX2_X2 U11624 ( .A(regBoiz_regfile_20__22_), .B(regBoiz_regfile_28__22_), 
        .S(net377166), .Z(n7747) );
  NAND2_X2 U11625 ( .A1(n7747), .A2(net367005), .ZN(n9856) );
  MUX2_X2 U11626 ( .A(regBoiz_regfile_17__22_), .B(regBoiz_regfile_25__22_), 
        .S(net369202), .Z(n7749) );
  MUX2_X2 U11627 ( .A(regBoiz_regfile_19__22_), .B(regBoiz_regfile_27__22_), 
        .S(net366899), .Z(n7748) );
  MUX2_X2 U11628 ( .A(n7749), .B(n7748), .S(net366977), .Z(n9853) );
  INV_X4 U11629 ( .A(n9853), .ZN(n7750) );
  NOR2_X4 U11630 ( .A1(n7750), .A2(n9854), .ZN(n7751) );
  NOR3_X4 U11631 ( .A1(n7753), .A2(n7752), .A3(n7751), .ZN(n7766) );
  MUX2_X2 U11632 ( .A(regBoiz_regfile_1__22_), .B(regBoiz_regfile_9__22_), .S(
        net366887), .Z(n7755) );
  MUX2_X2 U11633 ( .A(regBoiz_regfile_3__22_), .B(regBoiz_regfile_11__22_), 
        .S(net366887), .Z(n7754) );
  MUX2_X2 U11634 ( .A(n7755), .B(n7754), .S(net366973), .Z(n9851) );
  NAND2_X2 U11635 ( .A1(n9846), .A2(n9851), .ZN(n7765) );
  MUX2_X2 U11636 ( .A(regBoiz_regfile_16__22_), .B(regBoiz_regfile_24__22_), 
        .S(net377166), .Z(n7757) );
  MUX2_X2 U11637 ( .A(n7757), .B(n7756), .S(net366973), .Z(n9849) );
  INV_X4 U11638 ( .A(n9849), .ZN(n7758) );
  MUX2_X2 U11639 ( .A(regBoiz_regfile_21__22_), .B(regBoiz_regfile_29__22_), 
        .S(net377166), .Z(n7760) );
  MUX2_X2 U11640 ( .A(regBoiz_regfile_23__22_), .B(regBoiz_regfile_31__22_), 
        .S(net377166), .Z(n7759) );
  MUX2_X2 U11641 ( .A(n7760), .B(n7759), .S(net366973), .Z(n9861) );
  INV_X4 U11642 ( .A(n9861), .ZN(n7761) );
  NAND2_X2 U11643 ( .A1(n7944), .A2(net378321), .ZN(n9862) );
  OAI21_X4 U11644 ( .B1(n7761), .B2(n9862), .A(n9822), .ZN(n7762) );
  NOR2_X4 U11645 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  NAND2_X2 U11646 ( .A1(daddr[9]), .A2(n8157), .ZN(n9875) );
  INV_X4 U11647 ( .A(n9875), .ZN(n7767) );
  AOI21_X4 U11648 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n11112) );
  MUX2_X2 U11649 ( .A(regBoiz_regfile_1__23_), .B(regBoiz_regfile_5__23_), .S(
        regBoiz_N12), .Z(n7771) );
  MUX2_X2 U11650 ( .A(regBoiz_regfile_3__23_), .B(regBoiz_regfile_7__23_), .S(
        regBoiz_N12), .Z(n7770) );
  MUX2_X2 U11651 ( .A(n7771), .B(n7770), .S(net366973), .Z(n7775) );
  MUX2_X2 U11652 ( .A(regBoiz_regfile_17__23_), .B(regBoiz_regfile_21__23_), 
        .S(regBoiz_N12), .Z(n7773) );
  MUX2_X2 U11653 ( .A(regBoiz_regfile_9__23_), .B(regBoiz_regfile_13__23_), 
        .S(net366927), .Z(n7777) );
  MUX2_X2 U11654 ( .A(n7777), .B(n7776), .S(net366973), .Z(n7781) );
  MUX2_X2 U11655 ( .A(regBoiz_regfile_27__23_), .B(n6378), .S(regBoiz_N12), 
        .Z(n7778) );
  OAI21_X4 U11656 ( .B1(n7788), .B2(n7787), .A(net366999), .ZN(n7796) );
  NAND2_X2 U11657 ( .A1(regBoiz_regfile_14__23_), .A2(net375727), .ZN(n7789)
         );
  NAND2_X2 U11658 ( .A1(regBoiz_regfile_10__23_), .A2(net376330), .ZN(n7791)
         );
  OAI21_X4 U11659 ( .B1(n7794), .B2(n7793), .A(net366969), .ZN(n7795) );
  MUX2_X2 U11660 ( .A(regBoiz_regfile_16__23_), .B(regBoiz_regfile_24__23_), 
        .S(net366885), .Z(n7798) );
  MUX2_X2 U11661 ( .A(n7798), .B(n7797), .S(net366973), .Z(n7802) );
  MUX2_X2 U11662 ( .A(n7802), .B(n7801), .S(net366939), .Z(n9878) );
  MUX2_X2 U11663 ( .A(regBoiz_regfile_9__24_), .B(regBoiz_regfile_25__24_), 
        .S(n6788), .Z(n7807) );
  INV_X4 U11664 ( .A(n7807), .ZN(n7808) );
  INV_X4 U11665 ( .A(net365284), .ZN(net365293) );
  MUX2_X2 U11666 ( .A(regBoiz_regfile_15__24_), .B(regBoiz_regfile_31__24_), 
        .S(n6788), .Z(n7809) );
  INV_X4 U11667 ( .A(n7809), .ZN(n7810) );
  NAND2_X2 U11668 ( .A1(n7812), .A2(n7811), .ZN(n7864) );
  MUX2_X2 U11669 ( .A(regBoiz_regfile_11__24_), .B(regBoiz_regfile_27__24_), 
        .S(n6788), .Z(n7813) );
  INV_X4 U11670 ( .A(n7813), .ZN(n7814) );
  MUX2_X2 U11671 ( .A(regBoiz_regfile_13__24_), .B(regBoiz_regfile_29__24_), 
        .S(n6788), .Z(n7815) );
  INV_X4 U11672 ( .A(n7815), .ZN(n7816) );
  NAND2_X2 U11673 ( .A1(regBoiz_regfile_7__24_), .A2(n6795), .ZN(n7818) );
  NAND2_X2 U11674 ( .A1(regBoiz_regfile_23__24_), .A2(n6787), .ZN(n7817) );
  AOI21_X4 U11675 ( .B1(n7818), .B2(n7817), .A(net366951), .ZN(n7822) );
  NAND2_X2 U11676 ( .A1(regBoiz_regfile_3__24_), .A2(n6795), .ZN(n7820) );
  NAND2_X2 U11677 ( .A1(regBoiz_regfile_5__24_), .A2(n6795), .ZN(n7824) );
  NAND2_X2 U11678 ( .A1(regBoiz_regfile_21__24_), .A2(n6788), .ZN(n7823) );
  NAND2_X2 U11679 ( .A1(regBoiz_regfile_1__24_), .A2(n6795), .ZN(n7826) );
  NAND2_X2 U11680 ( .A1(regBoiz_regfile_17__24_), .A2(n6787), .ZN(n7825) );
  NAND4_X2 U11681 ( .A1(n7833), .A2(n7832), .A3(net367025), .A4(n7831), .ZN(
        n7863) );
  MUX2_X2 U11682 ( .A(regBoiz_regfile_4__24_), .B(regBoiz_regfile_12__24_), 
        .S(net366887), .Z(n7834) );
  INV_X4 U11683 ( .A(n7834), .ZN(n7835) );
  NOR2_X4 U11684 ( .A1(net366967), .A2(n6782), .ZN(n7841) );
  MUX2_X2 U11685 ( .A(regBoiz_regfile_6__24_), .B(regBoiz_regfile_14__24_), 
        .S(net366887), .Z(n7836) );
  INV_X4 U11686 ( .A(n7836), .ZN(n7837) );
  MUX2_X2 U11687 ( .A(regBoiz_regfile_2__24_), .B(regBoiz_regfile_10__24_), 
        .S(net376330), .Z(n7838) );
  INV_X4 U11688 ( .A(n7838), .ZN(n7839) );
  MUX2_X2 U11689 ( .A(regBoiz_regfile_0__24_), .B(regBoiz_regfile_8__24_), .S(
        net366887), .Z(n7840) );
  INV_X4 U11690 ( .A(n7840), .ZN(n7842) );
  NAND4_X2 U11691 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n7862)
         );
  MUX2_X2 U11692 ( .A(regBoiz_regfile_16__24_), .B(regBoiz_regfile_24__24_), 
        .S(net369202), .Z(n7847) );
  NAND2_X2 U11693 ( .A1(n6787), .A2(net367005), .ZN(n7850) );
  MUX2_X2 U11694 ( .A(regBoiz_regfile_20__24_), .B(regBoiz_regfile_28__24_), 
        .S(net376374), .Z(n7849) );
  INV_X4 U11695 ( .A(n7849), .ZN(n7852) );
  INV_X4 U11696 ( .A(n7850), .ZN(n7851) );
  MUX2_X2 U11697 ( .A(regBoiz_regfile_22__24_), .B(regBoiz_regfile_30__24_), 
        .S(net369202), .Z(n7853) );
  INV_X4 U11698 ( .A(n7853), .ZN(n7855) );
  NAND2_X2 U11699 ( .A1(n6787), .A2(net366987), .ZN(n7856) );
  INV_X4 U11700 ( .A(n7856), .ZN(n7854) );
  MUX2_X2 U11701 ( .A(regBoiz_regfile_18__24_), .B(regBoiz_regfile_26__24_), 
        .S(net369202), .Z(n7857) );
  NAND4_X2 U11702 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n5453), .ZN(n7861)
         );
  NAND2_X2 U11703 ( .A1(daddr[7]), .A2(net362342), .ZN(n9888) );
  OAI21_X4 U11704 ( .B1(n7865), .B2(net368548), .A(n9888), .ZN(n13536) );
  NAND2_X2 U11705 ( .A1(regBoiz_regfile_4__25_), .A2(n6795), .ZN(n7867) );
  NAND2_X2 U11706 ( .A1(regBoiz_regfile_20__25_), .A2(n6789), .ZN(n7866) );
  NAND2_X2 U11707 ( .A1(regBoiz_regfile_0__25_), .A2(n6795), .ZN(n7869) );
  NAND2_X2 U11708 ( .A1(regBoiz_regfile_16__25_), .A2(n6787), .ZN(n7868) );
  NAND2_X2 U11709 ( .A1(regBoiz_regfile_6__25_), .A2(n6795), .ZN(n7873) );
  NAND2_X2 U11710 ( .A1(regBoiz_regfile_22__25_), .A2(n6788), .ZN(n7872) );
  NAND2_X2 U11711 ( .A1(regBoiz_regfile_2__25_), .A2(n6795), .ZN(n7875) );
  NAND2_X2 U11712 ( .A1(regBoiz_regfile_18__25_), .A2(n6788), .ZN(n7874) );
  OAI21_X4 U11713 ( .B1(n7877), .B2(n7876), .A(net366969), .ZN(n7878) );
  NAND2_X2 U11714 ( .A1(regBoiz_regfile_12__25_), .A2(n6795), .ZN(n7881) );
  NAND2_X2 U11715 ( .A1(regBoiz_regfile_28__25_), .A2(n6787), .ZN(n7880) );
  NAND2_X2 U11716 ( .A1(regBoiz_regfile_8__25_), .A2(n6795), .ZN(n7883) );
  NAND2_X2 U11717 ( .A1(regBoiz_regfile_24__25_), .A2(n6787), .ZN(n7882) );
  OAI21_X4 U11718 ( .B1(n7885), .B2(n7884), .A(net367001), .ZN(n7893) );
  NAND2_X2 U11719 ( .A1(regBoiz_regfile_14__25_), .A2(n6795), .ZN(n7887) );
  NAND2_X2 U11720 ( .A1(regBoiz_regfile_30__25_), .A2(n6788), .ZN(n7886) );
  NAND2_X2 U11721 ( .A1(regBoiz_regfile_10__25_), .A2(n6795), .ZN(n7889) );
  NAND2_X2 U11722 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  MUX2_X2 U11723 ( .A(n7895), .B(n7894), .S(n5242), .Z(n7896) );
  NAND2_X2 U11724 ( .A1(regBoiz_regfile_5__25_), .A2(n6795), .ZN(n7898) );
  NAND2_X2 U11725 ( .A1(regBoiz_regfile_21__25_), .A2(n6788), .ZN(n7897) );
  NAND2_X2 U11726 ( .A1(regBoiz_regfile_1__25_), .A2(n6795), .ZN(n7900) );
  NAND2_X2 U11727 ( .A1(regBoiz_regfile_17__25_), .A2(n6788), .ZN(n7899) );
  OAI21_X4 U11728 ( .B1(n7902), .B2(n7901), .A(net366999), .ZN(n7910) );
  NAND2_X2 U11729 ( .A1(regBoiz_regfile_7__25_), .A2(n6795), .ZN(n7904) );
  NAND2_X2 U11730 ( .A1(regBoiz_regfile_23__25_), .A2(n6787), .ZN(n7903) );
  NAND2_X2 U11731 ( .A1(regBoiz_regfile_3__25_), .A2(n6794), .ZN(n7906) );
  NAND2_X2 U11732 ( .A1(regBoiz_regfile_19__25_), .A2(n6787), .ZN(n7905) );
  OAI21_X4 U11733 ( .B1(n7908), .B2(n7907), .A(net366969), .ZN(n7909) );
  NAND2_X2 U11734 ( .A1(n7910), .A2(n7909), .ZN(n7926) );
  NAND2_X2 U11735 ( .A1(regBoiz_regfile_13__25_), .A2(n6794), .ZN(n7912) );
  NAND2_X2 U11736 ( .A1(regBoiz_regfile_29__25_), .A2(n6788), .ZN(n7911) );
  NAND2_X2 U11737 ( .A1(regBoiz_regfile_9__25_), .A2(n6794), .ZN(n7914) );
  OAI21_X4 U11738 ( .B1(n7916), .B2(n7915), .A(net366999), .ZN(n7924) );
  NAND2_X2 U11739 ( .A1(regBoiz_regfile_15__25_), .A2(n6794), .ZN(n7918) );
  NAND2_X2 U11740 ( .A1(regBoiz_regfile_31__25_), .A2(n6787), .ZN(n7917) );
  NAND2_X2 U11741 ( .A1(regBoiz_regfile_11__25_), .A2(n6794), .ZN(n7920) );
  NAND2_X2 U11742 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  MUX2_X2 U11743 ( .A(n7926), .B(n7925), .S(n5242), .Z(n7927) );
  NAND2_X2 U11744 ( .A1(net367029), .A2(n7927), .ZN(n7928) );
  INV_X4 U11745 ( .A(n7928), .ZN(n9795) );
  NOR2_X4 U11746 ( .A1(n7929), .A2(n9795), .ZN(n7930) );
  NAND2_X2 U11747 ( .A1(daddr[6]), .A2(net362342), .ZN(n9792) );
  MUX2_X2 U11748 ( .A(regBoiz_regfile_16__26_), .B(regBoiz_regfile_24__26_), 
        .S(net369202), .Z(n7932) );
  MUX2_X2 U11749 ( .A(regBoiz_regfile_19__26_), .B(regBoiz_regfile_27__26_), 
        .S(net369202), .Z(n7940) );
  INV_X4 U11750 ( .A(n7933), .ZN(n7970) );
  MUX2_X2 U11751 ( .A(regBoiz_regfile_17__26_), .B(regBoiz_regfile_25__26_), 
        .S(net369202), .Z(n7939) );
  MUX2_X2 U11752 ( .A(regBoiz_regfile_22__26_), .B(regBoiz_regfile_30__26_), 
        .S(net369202), .Z(n7942) );
  NAND2_X2 U11753 ( .A1(n9855), .A2(net366987), .ZN(n7941) );
  MUX2_X2 U11754 ( .A(regBoiz_regfile_23__26_), .B(regBoiz_regfile_31__26_), 
        .S(net369202), .Z(n7946) );
  INV_X4 U11755 ( .A(n7943), .ZN(n7944) );
  NAND3_X4 U11756 ( .A1(net366919), .A2(net366965), .A3(n7944), .ZN(n7945) );
  NOR2_X4 U11757 ( .A1(n7947), .A2(n6531), .ZN(n7952) );
  MUX2_X2 U11758 ( .A(regBoiz_regfile_20__26_), .B(regBoiz_regfile_28__26_), 
        .S(net376331), .Z(n7949) );
  NAND2_X2 U11759 ( .A1(n9855), .A2(net367005), .ZN(n7948) );
  NAND3_X4 U11760 ( .A1(n5421), .A2(n7952), .A3(n7951), .ZN(n7953) );
  AOI211_X4 U11761 ( .C1(n5439), .C2(n8025), .A(n7953), .B(n7954), .ZN(n7962)
         );
  INV_X4 U11762 ( .A(n9848), .ZN(n9867) );
  MUX2_X2 U11763 ( .A(n5383), .B(n5589), .S(net376330), .Z(n7958) );
  MUX2_X2 U11764 ( .A(n5578), .B(n5341), .S(net369200), .Z(n7957) );
  MUX2_X2 U11765 ( .A(n7958), .B(n7957), .S(net366973), .Z(n7959) );
  NAND2_X2 U11766 ( .A1(n9867), .A2(net367045), .ZN(net365106) );
  INV_X4 U11767 ( .A(net365106), .ZN(net365093) );
  MUX2_X2 U11768 ( .A(regBoiz_regfile_4__26_), .B(regBoiz_regfile_12__26_), 
        .S(net376330), .Z(n7964) );
  NAND2_X2 U11769 ( .A1(net365093), .A2(n7965), .ZN(n7968) );
  NAND2_X2 U11770 ( .A1(n9846), .A2(net367045), .ZN(net363057) );
  MUX2_X2 U11771 ( .A(regBoiz_regfile_0__26_), .B(regBoiz_regfile_8__26_), .S(
        net376331), .Z(n7967) );
  MUX2_X2 U11772 ( .A(regBoiz_regfile_23__27_), .B(regBoiz_regfile_31__27_), 
        .S(net376374), .Z(n7974) );
  INV_X4 U11773 ( .A(n7976), .ZN(n7972) );
  NAND2_X2 U11774 ( .A1(n7972), .A2(net366987), .ZN(n7973) );
  MUX2_X2 U11775 ( .A(regBoiz_regfile_21__27_), .B(regBoiz_regfile_29__27_), 
        .S(net366887), .Z(n7977) );
  NOR2_X4 U11776 ( .A1(n7977), .A2(n5441), .ZN(n7978) );
  INV_X4 U11777 ( .A(n7978), .ZN(n7979) );
  MUX2_X2 U11778 ( .A(regBoiz_regfile_20__27_), .B(regBoiz_regfile_28__27_), 
        .S(net376374), .Z(n7981) );
  MUX2_X2 U11779 ( .A(regBoiz_regfile_22__27_), .B(regBoiz_regfile_30__27_), 
        .S(net377166), .Z(n7982) );
  INV_X4 U11780 ( .A(n7982), .ZN(n7984) );
  NAND2_X2 U11781 ( .A1(n5454), .A2(n7985), .ZN(n7986) );
  NOR2_X4 U11782 ( .A1(n7987), .A2(n7986), .ZN(net365030) );
  MUX2_X2 U11783 ( .A(n5336), .B(n5419), .S(net368770), .Z(n7988) );
  MUX2_X2 U11784 ( .A(regBoiz_regfile_17__27_), .B(regBoiz_regfile_25__27_), 
        .S(net376077), .Z(n7991) );
  MUX2_X2 U11785 ( .A(n5337), .B(n5423), .S(net366887), .Z(n7995) );
  MUX2_X2 U11786 ( .A(n5338), .B(n5424), .S(net375510), .Z(n7994) );
  MUX2_X2 U11787 ( .A(n5339), .B(n5425), .S(net366885), .Z(n7998) );
  MUX2_X2 U11788 ( .A(n5340), .B(n5426), .S(net375510), .Z(n7997) );
  MUX2_X2 U11789 ( .A(regBoiz_regfile_1__28_), .B(n6018), .S(n6370), .Z(n8001)
         );
  MUX2_X2 U11790 ( .A(n8001), .B(n8000), .S(net366987), .Z(n8002) );
  NOR2_X4 U11791 ( .A1(n8122), .A2(n8002), .ZN(n10476) );
  MUX2_X2 U11792 ( .A(regBoiz_regfile_5__28_), .B(regBoiz_regfile_21__28_), 
        .S(n6783), .Z(n8004) );
  MUX2_X2 U11793 ( .A(regBoiz_regfile_15__28_), .B(regBoiz_regfile_31__28_), 
        .S(n6788), .Z(n8006) );
  OAI21_X4 U11794 ( .B1(n8006), .B2(n8005), .A(net364906), .ZN(n8010) );
  MUX2_X2 U11795 ( .A(regBoiz_regfile_7__28_), .B(regBoiz_regfile_23__28_), 
        .S(n6783), .Z(n8008) );
  NOR3_X4 U11796 ( .A1(n8011), .A2(n8010), .A3(n8009), .ZN(n8024) );
  MUX2_X2 U11797 ( .A(regBoiz_regfile_11__28_), .B(regBoiz_regfile_27__28_), 
        .S(n6788), .Z(n8014) );
  NAND3_X4 U11798 ( .A1(net366947), .A2(n8012), .A3(net366965), .ZN(n8013) );
  NOR2_X4 U11799 ( .A1(n8014), .A2(n8013), .ZN(n8022) );
  MUX2_X2 U11800 ( .A(regBoiz_regfile_9__28_), .B(regBoiz_regfile_25__28_), 
        .S(n6783), .Z(n8017) );
  NOR2_X4 U11801 ( .A1(n8017), .A2(n8016), .ZN(n8021) );
  MUX2_X2 U11802 ( .A(regBoiz_regfile_13__28_), .B(regBoiz_regfile_29__28_), 
        .S(n6788), .Z(n8019) );
  NOR3_X4 U11803 ( .A1(n8022), .A2(n8021), .A3(n8020), .ZN(n8023) );
  INV_X4 U11804 ( .A(n8025), .ZN(n9850) );
  MUX2_X2 U11805 ( .A(n8027), .B(n8026), .S(net366977), .Z(n8032) );
  MUX2_X2 U11806 ( .A(regBoiz_regfile_12__28_), .B(regBoiz_regfile_28__28_), 
        .S(n6789), .Z(n8029) );
  MUX2_X2 U11807 ( .A(regBoiz_regfile_14__28_), .B(regBoiz_regfile_30__28_), 
        .S(n6796), .Z(n8028) );
  MUX2_X2 U11808 ( .A(regBoiz_regfile_4__28_), .B(regBoiz_regfile_20__28_), 
        .S(n6789), .Z(n8036) );
  MUX2_X2 U11809 ( .A(regBoiz_regfile_6__28_), .B(regBoiz_regfile_22__28_), 
        .S(n6783), .Z(n8035) );
  MUX2_X2 U11810 ( .A(n8036), .B(n8035), .S(net366987), .Z(n8037) );
  INV_X4 U11811 ( .A(n8039), .ZN(n8122) );
  MUX2_X2 U11812 ( .A(regBoiz_regfile_0__28_), .B(regBoiz_regfile_16__28_), 
        .S(n6783), .Z(n8041) );
  MUX2_X2 U11813 ( .A(regBoiz_regfile_1__29_), .B(regBoiz_regfile_9__29_), .S(
        net366887), .Z(n8045) );
  MUX2_X2 U11814 ( .A(regBoiz_regfile_3__29_), .B(n6031), .S(net375510), .Z(
        n8044) );
  MUX2_X2 U11815 ( .A(n8045), .B(n8044), .S(net366987), .Z(n10435) );
  MUX2_X2 U11816 ( .A(regBoiz_regfile_5__29_), .B(regBoiz_regfile_13__29_), 
        .S(net366887), .Z(n8046) );
  NAND2_X2 U11817 ( .A1(n8046), .A2(net367005), .ZN(n10433) );
  MUX2_X2 U11818 ( .A(regBoiz_regfile_7__29_), .B(regBoiz_regfile_15__29_), 
        .S(net366887), .Z(n8047) );
  NAND2_X2 U11819 ( .A1(net366987), .A2(n8047), .ZN(n10432) );
  NAND3_X2 U11820 ( .A1(n10433), .A2(n10432), .A3(net366919), .ZN(n8048) );
  NAND2_X2 U11821 ( .A1(n11053), .A2(n8048), .ZN(n8058) );
  MUX2_X2 U11822 ( .A(regBoiz_regfile_6__29_), .B(n6172), .S(net375642), .Z(
        net364971) );
  NAND2_X2 U11823 ( .A1(n6531), .A2(net364803), .ZN(n8053) );
  MUX2_X2 U11824 ( .A(regBoiz_regfile_17__29_), .B(regBoiz_regfile_25__29_), 
        .S(net366899), .Z(n8065) );
  MUX2_X2 U11825 ( .A(regBoiz_regfile_19__29_), .B(regBoiz_regfile_27__29_), 
        .S(net368782), .Z(n8064) );
  MUX2_X2 U11826 ( .A(regBoiz_regfile_16__29_), .B(regBoiz_regfile_24__29_), 
        .S(net377166), .Z(n8068) );
  MUX2_X2 U11827 ( .A(regBoiz_regfile_18__29_), .B(n6176), .S(net366885), .Z(
        n8067) );
  MUX2_X2 U11828 ( .A(regBoiz_regfile_20__29_), .B(regBoiz_regfile_28__29_), 
        .S(net368781), .Z(n8071) );
  MUX2_X2 U11829 ( .A(regBoiz_regfile_22__29_), .B(n6284), .S(n5171), .Z(n8070) );
  NAND3_X2 U11830 ( .A1(n10437), .A2(n10436), .A3(net367043), .ZN(n8073) );
  NAND2_X2 U11831 ( .A1(regBoiz_regfile_10__30_), .A2(n6794), .ZN(n8075) );
  NAND2_X2 U11832 ( .A1(regBoiz_regfile_30__30_), .A2(n6788), .ZN(n8077) );
  OAI211_X2 U11833 ( .C1(n6787), .C2(n5408), .A(net378321), .B(n8077), .ZN(
        n8083) );
  NAND2_X2 U11834 ( .A1(regBoiz_regfile_8__30_), .A2(n6794), .ZN(n8078) );
  NAND2_X2 U11835 ( .A1(regBoiz_regfile_28__30_), .A2(n6788), .ZN(n8080) );
  OAI211_X2 U11836 ( .C1(n6787), .C2(n5409), .A(net366919), .B(n8080), .ZN(
        n8081) );
  NOR3_X4 U11837 ( .A1(n8157), .A2(n8086), .A3(n8085), .ZN(n8087) );
  NOR2_X4 U11838 ( .A1(n8088), .A2(n8087), .ZN(net364870) );
  NAND2_X2 U11839 ( .A1(regBoiz_regfile_4__30_), .A2(n6794), .ZN(n8090) );
  NAND2_X2 U11840 ( .A1(regBoiz_regfile_20__30_), .A2(n6788), .ZN(n8089) );
  NAND2_X2 U11841 ( .A1(regBoiz_regfile_16__30_), .A2(n6788), .ZN(n8091) );
  NAND2_X2 U11842 ( .A1(regBoiz_regfile_6__30_), .A2(n6794), .ZN(n8096) );
  NAND2_X2 U11843 ( .A1(regBoiz_regfile_22__30_), .A2(n6788), .ZN(n8095) );
  NAND2_X2 U11844 ( .A1(regBoiz_regfile_18__30_), .A2(n6788), .ZN(n8097) );
  NAND2_X2 U11845 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  MUX2_X2 U11846 ( .A(regBoiz_regfile_5__30_), .B(regBoiz_regfile_21__30_), 
        .S(n6783), .Z(n8104) );
  MUX2_X2 U11847 ( .A(regBoiz_regfile_7__30_), .B(regBoiz_regfile_23__30_), 
        .S(n6788), .Z(n8105) );
  NOR3_X4 U11848 ( .A1(n8106), .A2(n8105), .A3(net366997), .ZN(net364899) );
  NAND2_X2 U11849 ( .A1(regBoiz_regfile_15__30_), .A2(n6794), .ZN(n8108) );
  NAND2_X2 U11850 ( .A1(regBoiz_regfile_31__30_), .A2(n6788), .ZN(n8107) );
  NAND2_X2 U11851 ( .A1(regBoiz_regfile_27__30_), .A2(n6788), .ZN(n8109) );
  NAND2_X2 U11852 ( .A1(regBoiz_regfile_13__30_), .A2(n6794), .ZN(n8114) );
  NAND2_X2 U11853 ( .A1(regBoiz_regfile_29__30_), .A2(n6788), .ZN(n8113) );
  NAND2_X2 U11854 ( .A1(regBoiz_regfile_9__30_), .A2(n6794), .ZN(n8116) );
  NAND2_X2 U11855 ( .A1(regBoiz_regfile_25__30_), .A2(n6788), .ZN(n8115) );
  MUX2_X2 U11856 ( .A(regBoiz_regfile_3__30_), .B(regBoiz_regfile_19__30_), 
        .S(n6783), .Z(n8121) );
  MUX2_X2 U11857 ( .A(regBoiz_regfile_1__30_), .B(regBoiz_regfile_17__30_), 
        .S(n6783), .Z(n8123) );
  NAND2_X2 U11858 ( .A1(regBoiz_regfile_25__31_), .A2(n6788), .ZN(n8127) );
  NAND2_X2 U11859 ( .A1(regBoiz_regfile_27__31_), .A2(n6788), .ZN(n8128) );
  OAI211_X2 U11860 ( .C1(n6787), .C2(n5570), .A(n8128), .B(net366951), .ZN(
        n8129) );
  OAI22_X2 U11861 ( .A1(n8130), .A2(n8150), .B1(n8129), .B2(n8152), .ZN(n8141)
         );
  NAND2_X2 U11862 ( .A1(regBoiz_regfile_19__31_), .A2(n6788), .ZN(n8131) );
  NAND2_X2 U11863 ( .A1(n8131), .A2(net366953), .ZN(n8132) );
  NOR3_X4 U11864 ( .A1(n8134), .A2(n8133), .A3(n8132), .ZN(n8140) );
  NAND2_X2 U11865 ( .A1(regBoiz_regfile_17__31_), .A2(n6788), .ZN(n8135) );
  NAND2_X2 U11866 ( .A1(n8135), .A2(net366953), .ZN(n8136) );
  NOR3_X4 U11867 ( .A1(n8138), .A2(n8137), .A3(n8136), .ZN(n8139) );
  NOR3_X4 U11868 ( .A1(n8141), .A2(n8140), .A3(n8139), .ZN(n8160) );
  NAND2_X2 U11869 ( .A1(regBoiz_regfile_21__31_), .A2(n6788), .ZN(n8143) );
  NAND2_X2 U11870 ( .A1(regBoiz_regfile_23__31_), .A2(n6788), .ZN(n8146) );
  NAND2_X2 U11871 ( .A1(n8149), .A2(n8148), .ZN(n8156) );
  NOR3_X4 U11872 ( .A1(n8156), .A2(n8155), .A3(n8154), .ZN(n8159) );
  NOR2_X4 U11873 ( .A1(n8157), .A2(net367041), .ZN(n8158) );
  NAND3_X4 U11874 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(net362281) );
  MUX2_X2 U11875 ( .A(regBoiz_regfile_16__31_), .B(regBoiz_regfile_24__31_), 
        .S(net369204), .Z(n8161) );
  INV_X4 U11876 ( .A(n8161), .ZN(n8164) );
  MUX2_X2 U11877 ( .A(regBoiz_regfile_18__31_), .B(regBoiz_regfile_26__31_), 
        .S(net377166), .Z(n8162) );
  MUX2_X2 U11878 ( .A(regBoiz_regfile_22__31_), .B(regBoiz_regfile_30__31_), 
        .S(net369204), .Z(n8165) );
  NAND2_X2 U11879 ( .A1(net366987), .A2(n8165), .ZN(n8168) );
  MUX2_X2 U11880 ( .A(regBoiz_regfile_20__31_), .B(regBoiz_regfile_28__31_), 
        .S(net368781), .Z(n8166) );
  NAND2_X2 U11881 ( .A1(n8166), .A2(net367005), .ZN(n8167) );
  NAND3_X2 U11882 ( .A1(n8168), .A2(n8167), .A3(net378321), .ZN(n8169) );
  AOI21_X4 U11883 ( .B1(n8171), .B2(net366949), .A(n8170), .ZN(n8183) );
  MUX2_X2 U11884 ( .A(n8173), .B(n8172), .S(net375527), .Z(n8174) );
  NAND2_X2 U11885 ( .A1(n9867), .A2(n8174), .ZN(n8179) );
  MUX2_X2 U11886 ( .A(regBoiz_regfile_0__31_), .B(regBoiz_regfile_8__31_), .S(
        n5248), .Z(n8176) );
  NAND2_X2 U11887 ( .A1(net364803), .A2(net367045), .ZN(n8180) );
  NAND2_X2 U11888 ( .A1(n6835), .A2(n6832), .ZN(n8190) );
  MUX2_X2 U11889 ( .A(regBoiz_regfile_24__27_), .B(regBoiz_regfile_25__27_), 
        .S(net369145), .Z(n8185) );
  MUX2_X2 U11890 ( .A(regBoiz_regfile_26__27_), .B(regBoiz_regfile_27__27_), 
        .S(net369162), .Z(n8184) );
  MUX2_X2 U11891 ( .A(n8185), .B(n8184), .S(n6799), .Z(n13001) );
  NAND2_X2 U11892 ( .A1(n8186), .A2(n13001), .ZN(n8196) );
  MUX2_X2 U11893 ( .A(regBoiz_regfile_20__27_), .B(regBoiz_regfile_21__27_), 
        .S(net369144), .Z(n8188) );
  MUX2_X2 U11894 ( .A(regBoiz_regfile_22__27_), .B(regBoiz_regfile_23__27_), 
        .S(net369163), .Z(n8187) );
  MUX2_X2 U11895 ( .A(n8188), .B(n8187), .S(n6809), .Z(n12998) );
  NAND2_X2 U11896 ( .A1(n8189), .A2(n12998), .ZN(n8195) );
  MUX2_X2 U11897 ( .A(regBoiz_regfile_28__27_), .B(regBoiz_regfile_29__27_), 
        .S(net369165), .Z(n8192) );
  MUX2_X2 U11898 ( .A(regBoiz_regfile_30__27_), .B(regBoiz_regfile_31__27_), 
        .S(net369236), .Z(n8191) );
  MUX2_X2 U11899 ( .A(n8192), .B(n8191), .S(n6806), .Z(n13000) );
  NOR2_X4 U11900 ( .A1(n6834), .A2(n6830), .ZN(n8220) );
  AOI21_X4 U11901 ( .B1(n8193), .B2(n13000), .A(n8220), .ZN(n8194) );
  MUX2_X2 U11902 ( .A(regBoiz_regfile_12__27_), .B(regBoiz_regfile_13__27_), 
        .S(net369236), .Z(n8198) );
  MUX2_X2 U11903 ( .A(n8198), .B(n8197), .S(n6806), .Z(n12994) );
  NAND2_X2 U11904 ( .A1(n8199), .A2(n12994), .ZN(n8207) );
  MUX2_X2 U11905 ( .A(regBoiz_regfile_16__27_), .B(regBoiz_regfile_17__27_), 
        .S(net369147), .Z(n8201) );
  MUX2_X2 U11906 ( .A(regBoiz_regfile_18__27_), .B(regBoiz_regfile_19__27_), 
        .S(net369144), .Z(n8200) );
  MUX2_X2 U11907 ( .A(n8201), .B(n8200), .S(n6807), .Z(n12999) );
  NAND2_X2 U11908 ( .A1(n8202), .A2(n12999), .ZN(n8206) );
  MUX2_X2 U11909 ( .A(regBoiz_regfile_8__27_), .B(regBoiz_regfile_9__27_), .S(
        net378318), .Z(n8203) );
  MUX2_X2 U11910 ( .A(n8203), .B(net364779), .S(n6807), .Z(n12995) );
  NAND2_X2 U11911 ( .A1(n8204), .A2(n12995), .ZN(n8205) );
  NAND3_X2 U11912 ( .A1(n8207), .A2(n8206), .A3(n8205), .ZN(n8225) );
  XOR2_X2 U11913 ( .A(n6799), .B(aluRw[1]), .Z(n8209) );
  XOR2_X2 U11914 ( .A(net369212), .B(aluRw[0]), .Z(n8208) );
  NOR2_X4 U11915 ( .A1(n8209), .A2(n8208), .ZN(n8214) );
  XNOR2_X2 U11916 ( .A(n6834), .B(aluRw[4]), .ZN(n8213) );
  XOR2_X2 U11917 ( .A(n6830), .B(aluRw[3]), .Z(n8211) );
  XOR2_X2 U11918 ( .A(n6821), .B(aluRw[2]), .Z(n8210) );
  NOR2_X4 U11919 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  NAND3_X4 U11920 ( .A1(n8214), .A2(n8213), .A3(n8212), .ZN(n12925) );
  INV_X4 U11921 ( .A(n6556), .ZN(n8834) );
  NAND3_X4 U11922 ( .A1(n12925), .A2(n12926), .A3(n8834), .ZN(n8708) );
  MUX2_X2 U11923 ( .A(regBoiz_regfile_0__27_), .B(regBoiz_regfile_1__27_), .S(
        net369166), .Z(n8216) );
  MUX2_X2 U11924 ( .A(n8216), .B(net364764), .S(n6807), .Z(n12993) );
  NAND2_X2 U11925 ( .A1(n8220), .A2(n6829), .ZN(n8217) );
  NOR2_X4 U11926 ( .A1(n12993), .A2(n8217), .ZN(n8223) );
  MUX2_X2 U11927 ( .A(regBoiz_regfile_4__27_), .B(regBoiz_regfile_5__27_), .S(
        net369164), .Z(n8219) );
  MUX2_X2 U11928 ( .A(regBoiz_regfile_6__27_), .B(regBoiz_regfile_7__27_), .S(
        net369165), .Z(n8218) );
  MUX2_X2 U11929 ( .A(n8219), .B(n8218), .S(n6807), .Z(n12992) );
  NAND2_X2 U11930 ( .A1(n6823), .A2(n8220), .ZN(n8221) );
  NOR2_X4 U11931 ( .A1(n12992), .A2(n8221), .ZN(n8222) );
  OAI21_X4 U11932 ( .B1(n8226), .B2(n8225), .A(n8224), .ZN(n8229) );
  INV_X4 U11933 ( .A(n12925), .ZN(n12927) );
  NAND2_X2 U11934 ( .A1(n12927), .A2(n8834), .ZN(n8227) );
  NAND2_X2 U11935 ( .A1(daddr[4]), .A2(n6547), .ZN(n8228) );
  MUX2_X2 U11936 ( .A(regBoiz_regfile_0__28_), .B(regBoiz_regfile_1__28_), .S(
        net369164), .Z(n8232) );
  MUX2_X2 U11937 ( .A(regBoiz_regfile_2__28_), .B(regBoiz_regfile_3__28_), .S(
        net369162), .Z(n8231) );
  MUX2_X2 U11938 ( .A(n8232), .B(n8231), .S(n6807), .Z(n8236) );
  MUX2_X2 U11939 ( .A(regBoiz_regfile_4__28_), .B(regBoiz_regfile_5__28_), .S(
        net369166), .Z(n8234) );
  MUX2_X2 U11940 ( .A(regBoiz_regfile_6__28_), .B(regBoiz_regfile_7__28_), .S(
        net369145), .Z(n8233) );
  MUX2_X2 U11941 ( .A(n8234), .B(n8233), .S(n6807), .Z(n8235) );
  MUX2_X2 U11942 ( .A(n8236), .B(n8235), .S(n6823), .Z(n8244) );
  MUX2_X2 U11943 ( .A(regBoiz_regfile_8__28_), .B(regBoiz_regfile_9__28_), .S(
        net369165), .Z(n8238) );
  MUX2_X2 U11944 ( .A(regBoiz_regfile_10__28_), .B(regBoiz_regfile_11__28_), 
        .S(net369147), .Z(n8237) );
  MUX2_X2 U11945 ( .A(n8238), .B(n8237), .S(n6807), .Z(n8242) );
  MUX2_X2 U11946 ( .A(regBoiz_regfile_12__28_), .B(regBoiz_regfile_13__28_), 
        .S(net369144), .Z(n8240) );
  MUX2_X2 U11947 ( .A(regBoiz_regfile_14__28_), .B(regBoiz_regfile_15__28_), 
        .S(net369212), .Z(n8239) );
  MUX2_X2 U11948 ( .A(n8240), .B(n8239), .S(n6807), .Z(n8241) );
  MUX2_X2 U11949 ( .A(n8242), .B(n8241), .S(n6822), .Z(n8243) );
  MUX2_X2 U11950 ( .A(n8244), .B(n8243), .S(n6832), .Z(n8260) );
  MUX2_X2 U11951 ( .A(regBoiz_regfile_16__28_), .B(regBoiz_regfile_17__28_), 
        .S(net369164), .Z(n8246) );
  MUX2_X2 U11952 ( .A(regBoiz_regfile_18__28_), .B(regBoiz_regfile_19__28_), 
        .S(net369144), .Z(n8245) );
  MUX2_X2 U11953 ( .A(n8246), .B(n8245), .S(n6807), .Z(n8250) );
  MUX2_X2 U11954 ( .A(regBoiz_regfile_20__28_), .B(regBoiz_regfile_21__28_), 
        .S(net369165), .Z(n8248) );
  MUX2_X2 U11955 ( .A(regBoiz_regfile_22__28_), .B(regBoiz_regfile_23__28_), 
        .S(net369154), .Z(n8247) );
  MUX2_X2 U11956 ( .A(n8248), .B(n8247), .S(n6807), .Z(n8249) );
  MUX2_X2 U11957 ( .A(n8250), .B(n8249), .S(n6825), .Z(n8258) );
  MUX2_X2 U11958 ( .A(regBoiz_regfile_24__28_), .B(regBoiz_regfile_25__28_), 
        .S(net369145), .Z(n8252) );
  MUX2_X2 U11959 ( .A(regBoiz_regfile_26__28_), .B(regBoiz_regfile_27__28_), 
        .S(net369155), .Z(n8251) );
  MUX2_X2 U11960 ( .A(n8252), .B(n8251), .S(n6807), .Z(n8256) );
  MUX2_X2 U11961 ( .A(regBoiz_regfile_28__28_), .B(regBoiz_regfile_29__28_), 
        .S(net369156), .Z(n8254) );
  MUX2_X2 U11962 ( .A(regBoiz_regfile_30__28_), .B(regBoiz_regfile_31__28_), 
        .S(net369147), .Z(n8253) );
  MUX2_X2 U11963 ( .A(n8254), .B(n8253), .S(n6807), .Z(n8255) );
  MUX2_X2 U11964 ( .A(n8256), .B(n8255), .S(n6822), .Z(n8257) );
  MUX2_X2 U11965 ( .A(n8258), .B(n8257), .S(n6832), .Z(n8259) );
  MUX2_X2 U11966 ( .A(n8260), .B(n8259), .S(n6835), .Z(n13243) );
  NAND2_X2 U11967 ( .A1(n9718), .A2(n13243), .ZN(n8261) );
  NAND2_X2 U11968 ( .A1(daddr[3]), .A2(n6547), .ZN(n8698) );
  NAND2_X2 U11969 ( .A1(aluBoi_imm32w_2_), .A2(n6556), .ZN(n8294) );
  MUX2_X2 U11970 ( .A(regBoiz_regfile_0__29_), .B(regBoiz_regfile_1__29_), .S(
        net369162), .Z(n8263) );
  MUX2_X2 U11971 ( .A(regBoiz_regfile_2__29_), .B(regBoiz_regfile_3__29_), .S(
        net369162), .Z(n8262) );
  MUX2_X2 U11972 ( .A(n8263), .B(n8262), .S(n6801), .Z(n8267) );
  MUX2_X2 U11973 ( .A(regBoiz_regfile_4__29_), .B(regBoiz_regfile_5__29_), .S(
        net369147), .Z(n8265) );
  MUX2_X2 U11974 ( .A(n8265), .B(n8264), .S(n6802), .Z(n8266) );
  MUX2_X2 U11975 ( .A(n8267), .B(n8266), .S(n6823), .Z(n8275) );
  MUX2_X2 U11976 ( .A(regBoiz_regfile_8__29_), .B(regBoiz_regfile_9__29_), .S(
        net369242), .Z(n8269) );
  MUX2_X2 U11977 ( .A(regBoiz_regfile_10__29_), .B(regBoiz_regfile_11__29_), 
        .S(net369156), .Z(n8268) );
  MUX2_X2 U11978 ( .A(n8269), .B(n8268), .S(n6802), .Z(n8273) );
  MUX2_X2 U11979 ( .A(regBoiz_regfile_12__29_), .B(regBoiz_regfile_13__29_), 
        .S(net369222), .Z(n8271) );
  MUX2_X2 U11980 ( .A(regBoiz_regfile_14__29_), .B(regBoiz_regfile_15__29_), 
        .S(net377337), .Z(n8270) );
  MUX2_X2 U11981 ( .A(n8271), .B(n8270), .S(n6806), .Z(n8272) );
  MUX2_X2 U11982 ( .A(n8273), .B(n8272), .S(n6825), .Z(n8274) );
  MUX2_X2 U11983 ( .A(n8275), .B(n8274), .S(n6832), .Z(n8291) );
  MUX2_X2 U11984 ( .A(regBoiz_regfile_16__29_), .B(regBoiz_regfile_17__29_), 
        .S(net369145), .Z(n8277) );
  MUX2_X2 U11985 ( .A(regBoiz_regfile_18__29_), .B(regBoiz_regfile_19__29_), 
        .S(net369242), .Z(n8276) );
  MUX2_X2 U11986 ( .A(n8277), .B(n8276), .S(n6801), .Z(n8281) );
  MUX2_X2 U11987 ( .A(regBoiz_regfile_20__29_), .B(regBoiz_regfile_21__29_), 
        .S(net369144), .Z(n8279) );
  MUX2_X2 U11988 ( .A(regBoiz_regfile_22__29_), .B(regBoiz_regfile_23__29_), 
        .S(net369145), .Z(n8278) );
  MUX2_X2 U11989 ( .A(n8279), .B(n8278), .S(n6806), .Z(n8280) );
  MUX2_X2 U11990 ( .A(n8281), .B(n8280), .S(n6826), .Z(n8289) );
  MUX2_X2 U11991 ( .A(regBoiz_regfile_24__29_), .B(regBoiz_regfile_25__29_), 
        .S(net369234), .Z(n8283) );
  MUX2_X2 U11992 ( .A(regBoiz_regfile_26__29_), .B(regBoiz_regfile_27__29_), 
        .S(net369166), .Z(n8282) );
  MUX2_X2 U11993 ( .A(n8283), .B(n8282), .S(n6806), .Z(n8287) );
  MUX2_X2 U11994 ( .A(regBoiz_regfile_28__29_), .B(regBoiz_regfile_29__29_), 
        .S(net369147), .Z(n8285) );
  MUX2_X2 U11995 ( .A(regBoiz_regfile_30__29_), .B(regBoiz_regfile_31__29_), 
        .S(net369166), .Z(n8284) );
  MUX2_X2 U11996 ( .A(n8285), .B(n8284), .S(n6811), .Z(n8286) );
  MUX2_X2 U11997 ( .A(n8287), .B(n8286), .S(n6826), .Z(n8288) );
  MUX2_X2 U11998 ( .A(n8289), .B(n8288), .S(n6832), .Z(n8290) );
  MUX2_X2 U11999 ( .A(n8291), .B(n8290), .S(n6835), .Z(n13255) );
  NAND2_X2 U12000 ( .A1(n9718), .A2(n13255), .ZN(n8293) );
  NAND2_X2 U12001 ( .A1(daddr[2]), .A2(n6547), .ZN(n8292) );
  MUX2_X2 U12002 ( .A(regBoiz_regfile_0__30_), .B(regBoiz_regfile_1__30_), .S(
        net369218), .Z(n8296) );
  MUX2_X2 U12003 ( .A(regBoiz_regfile_2__30_), .B(regBoiz_regfile_3__30_), .S(
        net369154), .Z(n8295) );
  MUX2_X2 U12004 ( .A(n8296), .B(n8295), .S(n6806), .Z(n8300) );
  MUX2_X2 U12005 ( .A(regBoiz_regfile_4__30_), .B(regBoiz_regfile_5__30_), .S(
        net369218), .Z(n8298) );
  MUX2_X2 U12006 ( .A(regBoiz_regfile_6__30_), .B(regBoiz_regfile_7__30_), .S(
        net369218), .Z(n8297) );
  MUX2_X2 U12007 ( .A(n8298), .B(n8297), .S(n6809), .Z(n8299) );
  MUX2_X2 U12008 ( .A(n8300), .B(n8299), .S(n6826), .Z(n8308) );
  MUX2_X2 U12009 ( .A(regBoiz_regfile_8__30_), .B(regBoiz_regfile_9__30_), .S(
        net369155), .Z(n8302) );
  MUX2_X2 U12010 ( .A(regBoiz_regfile_10__30_), .B(regBoiz_regfile_11__30_), 
        .S(net369154), .Z(n8301) );
  MUX2_X2 U12011 ( .A(n8302), .B(n8301), .S(n6809), .Z(n8306) );
  MUX2_X2 U12012 ( .A(regBoiz_regfile_12__30_), .B(regBoiz_regfile_13__30_), 
        .S(net369155), .Z(n8304) );
  MUX2_X2 U12013 ( .A(regBoiz_regfile_14__30_), .B(regBoiz_regfile_15__30_), 
        .S(net369161), .Z(n8303) );
  MUX2_X2 U12014 ( .A(n8304), .B(n8303), .S(n6810), .Z(n8305) );
  MUX2_X2 U12015 ( .A(n8306), .B(n8305), .S(n6826), .Z(n8307) );
  MUX2_X2 U12016 ( .A(n8308), .B(n8307), .S(n6831), .Z(n8324) );
  MUX2_X2 U12017 ( .A(regBoiz_regfile_16__30_), .B(regBoiz_regfile_17__30_), 
        .S(net369144), .Z(n8310) );
  MUX2_X2 U12018 ( .A(regBoiz_regfile_18__30_), .B(regBoiz_regfile_19__30_), 
        .S(net369242), .Z(n8309) );
  MUX2_X2 U12019 ( .A(regBoiz_regfile_20__30_), .B(regBoiz_regfile_21__30_), 
        .S(net369147), .Z(n8312) );
  MUX2_X2 U12020 ( .A(regBoiz_regfile_22__30_), .B(regBoiz_regfile_23__30_), 
        .S(net369164), .Z(n8311) );
  MUX2_X2 U12021 ( .A(n8314), .B(n8313), .S(n6826), .Z(n8322) );
  MUX2_X2 U12022 ( .A(regBoiz_regfile_26__30_), .B(regBoiz_regfile_27__30_), 
        .S(net369162), .Z(n8315) );
  MUX2_X2 U12023 ( .A(n8316), .B(n8315), .S(n6808), .Z(n8320) );
  MUX2_X2 U12024 ( .A(regBoiz_regfile_28__30_), .B(regBoiz_regfile_29__30_), 
        .S(net369163), .Z(n8318) );
  MUX2_X2 U12025 ( .A(regBoiz_regfile_30__30_), .B(regBoiz_regfile_31__30_), 
        .S(n5770), .Z(n8317) );
  MUX2_X2 U12026 ( .A(n8318), .B(n8317), .S(n6808), .Z(n8319) );
  MUX2_X2 U12027 ( .A(n8322), .B(n8321), .S(n6832), .Z(n8323) );
  MUX2_X2 U12028 ( .A(n8324), .B(n8323), .S(n6835), .Z(n13266) );
  NAND2_X2 U12029 ( .A1(daddr[1]), .A2(n6547), .ZN(n8705) );
  MUX2_X2 U12030 ( .A(regBoiz_regfile_0__31_), .B(regBoiz_regfile_1__31_), .S(
        net377338), .Z(n8326) );
  MUX2_X2 U12031 ( .A(regBoiz_regfile_2__31_), .B(regBoiz_regfile_3__31_), .S(
        net369166), .Z(n8325) );
  MUX2_X2 U12032 ( .A(n8326), .B(n8325), .S(n6808), .Z(n8330) );
  MUX2_X2 U12033 ( .A(regBoiz_regfile_4__31_), .B(regBoiz_regfile_5__31_), .S(
        net369165), .Z(n8328) );
  MUX2_X2 U12034 ( .A(regBoiz_regfile_6__31_), .B(regBoiz_regfile_7__31_), .S(
        net369165), .Z(n8327) );
  MUX2_X2 U12035 ( .A(n8328), .B(n8327), .S(n6808), .Z(n8329) );
  MUX2_X2 U12036 ( .A(n8330), .B(n8329), .S(n6826), .Z(n8338) );
  MUX2_X2 U12037 ( .A(regBoiz_regfile_8__31_), .B(regBoiz_regfile_9__31_), .S(
        net369161), .Z(n8332) );
  MUX2_X2 U12038 ( .A(n8332), .B(n8331), .S(n6808), .Z(n8336) );
  MUX2_X2 U12039 ( .A(regBoiz_regfile_12__31_), .B(regBoiz_regfile_13__31_), 
        .S(net369161), .Z(n8334) );
  MUX2_X2 U12040 ( .A(regBoiz_regfile_14__31_), .B(regBoiz_regfile_15__31_), 
        .S(net369165), .Z(n8333) );
  MUX2_X2 U12041 ( .A(n8334), .B(n8333), .S(n6808), .Z(n8335) );
  MUX2_X2 U12042 ( .A(n8336), .B(n8335), .S(n6826), .Z(n8337) );
  MUX2_X2 U12043 ( .A(n8338), .B(n8337), .S(n6831), .Z(n8354) );
  MUX2_X2 U12044 ( .A(regBoiz_regfile_16__31_), .B(regBoiz_regfile_17__31_), 
        .S(net369155), .Z(n8340) );
  MUX2_X2 U12045 ( .A(regBoiz_regfile_18__31_), .B(regBoiz_regfile_19__31_), 
        .S(net369156), .Z(n8339) );
  MUX2_X2 U12046 ( .A(n8340), .B(n8339), .S(n6808), .Z(n8344) );
  MUX2_X2 U12047 ( .A(regBoiz_regfile_20__31_), .B(regBoiz_regfile_21__31_), 
        .S(net369155), .Z(n8342) );
  MUX2_X2 U12048 ( .A(regBoiz_regfile_22__31_), .B(regBoiz_regfile_23__31_), 
        .S(net369156), .Z(n8341) );
  MUX2_X2 U12049 ( .A(n8342), .B(n8341), .S(n6808), .Z(n8343) );
  MUX2_X2 U12050 ( .A(n8344), .B(n8343), .S(n6826), .Z(n8352) );
  MUX2_X2 U12051 ( .A(regBoiz_regfile_24__31_), .B(regBoiz_regfile_25__31_), 
        .S(net369166), .Z(n8346) );
  MUX2_X2 U12052 ( .A(regBoiz_regfile_26__31_), .B(regBoiz_regfile_27__31_), 
        .S(net369166), .Z(n8345) );
  MUX2_X2 U12053 ( .A(n8346), .B(n8345), .S(n6808), .Z(n8350) );
  MUX2_X2 U12054 ( .A(regBoiz_regfile_28__31_), .B(regBoiz_regfile_29__31_), 
        .S(net369214), .Z(n8348) );
  MUX2_X2 U12055 ( .A(n8354), .B(n8353), .S(n6835), .Z(n13277) );
  NAND2_X2 U12056 ( .A1(n9718), .A2(n13277), .ZN(n8355) );
  NAND2_X2 U12057 ( .A1(daddr[0]), .A2(n6547), .ZN(n8710) );
  NAND2_X2 U12058 ( .A1(idOut_24_), .A2(n5314), .ZN(n9189) );
  INV_X4 U12059 ( .A(n9189), .ZN(n9196) );
  INV_X4 U12060 ( .A(aluBoi_aluBoi_shft_sllout[9]), .ZN(n8362) );
  INV_X4 U12061 ( .A(aluBoi_aluBoi_shft_sllout[17]), .ZN(n8361) );
  INV_X4 U12062 ( .A(aluBoi_aluBoi_shft_sllout[16]), .ZN(n8360) );
  NAND4_X2 U12063 ( .A1(n8363), .A2(n8362), .A3(n8361), .A4(n8360), .ZN(n8364)
         );
  NAND2_X2 U12064 ( .A1(n8366), .A2(n8365), .ZN(n8382) );
  INV_X4 U12065 ( .A(aluBoi_aluBoi_shft_sraout[5]), .ZN(n8368) );
  INV_X4 U12066 ( .A(aluBoi_aluBoi_shft_sraout[0]), .ZN(n8372) );
  INV_X4 U12067 ( .A(aluBoi_aluBoi_shft_sraout[1]), .ZN(n8371) );
  INV_X4 U12068 ( .A(aluBoi_aluBoi_shft_sraout[2]), .ZN(n8370) );
  INV_X4 U12069 ( .A(aluBoi_aluBoi_shft_sraout[9]), .ZN(n8376) );
  NAND2_X2 U12070 ( .A1(idOut_22_), .A2(n9196), .ZN(n9766) );
  NAND2_X2 U12071 ( .A1(idOut_23_), .A2(n5314), .ZN(n9188) );
  INV_X4 U12072 ( .A(n13222), .ZN(n13220) );
  NAND2_X2 U12073 ( .A1(aluBoi_imm32w_14_), .A2(n6556), .ZN(n8415) );
  MUX2_X2 U12074 ( .A(regBoiz_regfile_0__17_), .B(regBoiz_regfile_1__17_), .S(
        net369244), .Z(n8384) );
  MUX2_X2 U12075 ( .A(regBoiz_regfile_2__17_), .B(regBoiz_regfile_3__17_), .S(
        net369214), .Z(n8383) );
  MUX2_X2 U12076 ( .A(n8384), .B(n8383), .S(n6801), .Z(n8388) );
  MUX2_X2 U12077 ( .A(regBoiz_regfile_4__17_), .B(regBoiz_regfile_5__17_), .S(
        net369156), .Z(n8386) );
  MUX2_X2 U12078 ( .A(regBoiz_regfile_6__17_), .B(regBoiz_regfile_7__17_), .S(
        net369228), .Z(n8385) );
  MUX2_X2 U12079 ( .A(n8386), .B(n8385), .S(n6804), .Z(n8387) );
  MUX2_X2 U12080 ( .A(n8388), .B(n8387), .S(n6826), .Z(n8396) );
  MUX2_X2 U12081 ( .A(regBoiz_regfile_8__17_), .B(regBoiz_regfile_9__17_), .S(
        net369157), .Z(n8390) );
  MUX2_X2 U12082 ( .A(regBoiz_regfile_10__17_), .B(regBoiz_regfile_11__17_), 
        .S(net369244), .Z(n8389) );
  MUX2_X2 U12083 ( .A(n8390), .B(n8389), .S(n6802), .Z(n8394) );
  MUX2_X2 U12084 ( .A(regBoiz_regfile_12__17_), .B(regBoiz_regfile_13__17_), 
        .S(net377338), .Z(n8392) );
  MUX2_X2 U12085 ( .A(regBoiz_regfile_14__17_), .B(regBoiz_regfile_15__17_), 
        .S(net369242), .Z(n8391) );
  MUX2_X2 U12086 ( .A(n8392), .B(n8391), .S(n6804), .Z(n8393) );
  MUX2_X2 U12087 ( .A(n8394), .B(n8393), .S(n6826), .Z(n8395) );
  MUX2_X2 U12088 ( .A(n8396), .B(n8395), .S(n6831), .Z(n8412) );
  MUX2_X2 U12089 ( .A(regBoiz_regfile_16__17_), .B(regBoiz_regfile_17__17_), 
        .S(net369165), .Z(n8398) );
  MUX2_X2 U12090 ( .A(regBoiz_regfile_18__17_), .B(regBoiz_regfile_19__17_), 
        .S(net369144), .Z(n8397) );
  MUX2_X2 U12091 ( .A(n8398), .B(n8397), .S(n6801), .Z(n8402) );
  MUX2_X2 U12092 ( .A(regBoiz_regfile_20__17_), .B(regBoiz_regfile_21__17_), 
        .S(net369161), .Z(n8400) );
  MUX2_X2 U12093 ( .A(regBoiz_regfile_22__17_), .B(regBoiz_regfile_23__17_), 
        .S(net369147), .Z(n8399) );
  MUX2_X2 U12094 ( .A(n8400), .B(n8399), .S(n6804), .Z(n8401) );
  MUX2_X2 U12095 ( .A(n8402), .B(n8401), .S(n6826), .Z(n8410) );
  MUX2_X2 U12096 ( .A(regBoiz_regfile_24__17_), .B(regBoiz_regfile_25__17_), 
        .S(net369145), .Z(n8404) );
  MUX2_X2 U12097 ( .A(regBoiz_regfile_26__17_), .B(regBoiz_regfile_27__17_), 
        .S(net369154), .Z(n8403) );
  MUX2_X2 U12098 ( .A(n8404), .B(n8403), .S(n6802), .Z(n8408) );
  MUX2_X2 U12099 ( .A(regBoiz_regfile_28__17_), .B(regBoiz_regfile_29__17_), 
        .S(net369155), .Z(n8406) );
  MUX2_X2 U12100 ( .A(regBoiz_regfile_30__17_), .B(regBoiz_regfile_31__17_), 
        .S(net377338), .Z(n8405) );
  MUX2_X2 U12101 ( .A(n8406), .B(n8405), .S(n6804), .Z(n8407) );
  MUX2_X2 U12102 ( .A(n8408), .B(n8407), .S(n6826), .Z(n8409) );
  MUX2_X2 U12103 ( .A(n8410), .B(n8409), .S(n6831), .Z(n8411) );
  MUX2_X2 U12104 ( .A(n8412), .B(n8411), .S(n6835), .Z(n12950) );
  NAND2_X2 U12105 ( .A1(n9718), .A2(n12950), .ZN(n8414) );
  NAND2_X2 U12106 ( .A1(daddr[14]), .A2(n6547), .ZN(n8413) );
  INV_X4 U12107 ( .A(n10418), .ZN(n9671) );
  XNOR2_X2 U12108 ( .A(n6565), .B(n9671), .ZN(n8767) );
  INV_X4 U12109 ( .A(n8935), .ZN(n9474) );
  NAND2_X2 U12110 ( .A1(aluBoi_imm32w_13_), .A2(n6556), .ZN(n8448) );
  MUX2_X2 U12111 ( .A(regBoiz_regfile_0__18_), .B(regBoiz_regfile_1__18_), .S(
        net369220), .Z(n8417) );
  MUX2_X2 U12112 ( .A(regBoiz_regfile_2__18_), .B(regBoiz_regfile_3__18_), .S(
        net369236), .Z(n8416) );
  MUX2_X2 U12113 ( .A(n8417), .B(n8416), .S(n6802), .Z(n8421) );
  MUX2_X2 U12114 ( .A(regBoiz_regfile_4__18_), .B(regBoiz_regfile_5__18_), .S(
        net369147), .Z(n8419) );
  MUX2_X2 U12115 ( .A(regBoiz_regfile_6__18_), .B(regBoiz_regfile_7__18_), .S(
        net369163), .Z(n8418) );
  MUX2_X2 U12116 ( .A(n8419), .B(n8418), .S(n6801), .Z(n8420) );
  MUX2_X2 U12117 ( .A(n8421), .B(n8420), .S(n6826), .Z(n8429) );
  MUX2_X2 U12118 ( .A(regBoiz_regfile_8__18_), .B(regBoiz_regfile_9__18_), .S(
        net369244), .Z(n8423) );
  MUX2_X2 U12119 ( .A(regBoiz_regfile_10__18_), .B(regBoiz_regfile_11__18_), 
        .S(net369165), .Z(n8422) );
  MUX2_X2 U12120 ( .A(n8423), .B(n8422), .S(n6804), .Z(n8427) );
  MUX2_X2 U12121 ( .A(regBoiz_regfile_12__18_), .B(regBoiz_regfile_13__18_), 
        .S(net369162), .Z(n8425) );
  MUX2_X2 U12122 ( .A(regBoiz_regfile_14__18_), .B(regBoiz_regfile_15__18_), 
        .S(net369161), .Z(n8424) );
  MUX2_X2 U12123 ( .A(n8425), .B(n8424), .S(n6802), .Z(n8426) );
  MUX2_X2 U12124 ( .A(n8427), .B(n8426), .S(n6826), .Z(n8428) );
  MUX2_X2 U12125 ( .A(n8429), .B(n8428), .S(n6831), .Z(n8445) );
  MUX2_X2 U12126 ( .A(regBoiz_regfile_16__18_), .B(regBoiz_regfile_17__18_), 
        .S(net378318), .Z(n8431) );
  MUX2_X2 U12127 ( .A(regBoiz_regfile_18__18_), .B(regBoiz_regfile_19__18_), 
        .S(net369214), .Z(n8430) );
  MUX2_X2 U12128 ( .A(n8431), .B(n8430), .S(n6804), .Z(n8435) );
  MUX2_X2 U12129 ( .A(regBoiz_regfile_20__18_), .B(regBoiz_regfile_21__18_), 
        .S(net369157), .Z(n8433) );
  MUX2_X2 U12130 ( .A(regBoiz_regfile_22__18_), .B(regBoiz_regfile_23__18_), 
        .S(net369166), .Z(n8432) );
  MUX2_X2 U12131 ( .A(n8433), .B(n8432), .S(n6804), .Z(n8434) );
  MUX2_X2 U12132 ( .A(n8435), .B(n8434), .S(n6825), .Z(n8443) );
  MUX2_X2 U12133 ( .A(regBoiz_regfile_24__18_), .B(regBoiz_regfile_25__18_), 
        .S(net369166), .Z(n8437) );
  MUX2_X2 U12134 ( .A(regBoiz_regfile_26__18_), .B(regBoiz_regfile_27__18_), 
        .S(net369214), .Z(n8436) );
  MUX2_X2 U12135 ( .A(n8437), .B(n8436), .S(n6804), .Z(n8441) );
  MUX2_X2 U12136 ( .A(regBoiz_regfile_28__18_), .B(regBoiz_regfile_29__18_), 
        .S(net369163), .Z(n8439) );
  MUX2_X2 U12137 ( .A(regBoiz_regfile_30__18_), .B(regBoiz_regfile_31__18_), 
        .S(net369164), .Z(n8438) );
  MUX2_X2 U12138 ( .A(n8439), .B(n8438), .S(n6804), .Z(n8440) );
  MUX2_X2 U12139 ( .A(n8441), .B(n8440), .S(n6825), .Z(n8442) );
  MUX2_X2 U12140 ( .A(n8443), .B(n8442), .S(n6831), .Z(n8444) );
  MUX2_X2 U12141 ( .A(n8445), .B(n8444), .S(n6835), .Z(n13055) );
  NAND2_X2 U12142 ( .A1(n9718), .A2(n13055), .ZN(n8447) );
  NAND2_X2 U12143 ( .A1(daddr[13]), .A2(n6547), .ZN(n8446) );
  INV_X4 U12144 ( .A(n10419), .ZN(n9661) );
  XNOR2_X2 U12145 ( .A(n6565), .B(n9661), .ZN(n8449) );
  INV_X4 U12146 ( .A(n8449), .ZN(n8450) );
  NAND2_X2 U12147 ( .A1(aluBoi_imm32w_10_), .A2(n6556), .ZN(n8483) );
  MUX2_X2 U12148 ( .A(regBoiz_regfile_0__21_), .B(regBoiz_regfile_1__21_), .S(
        net369226), .Z(n8452) );
  MUX2_X2 U12149 ( .A(regBoiz_regfile_2__21_), .B(regBoiz_regfile_3__21_), .S(
        net369144), .Z(n8451) );
  MUX2_X2 U12150 ( .A(n8452), .B(n8451), .S(n6801), .Z(n8456) );
  MUX2_X2 U12151 ( .A(regBoiz_regfile_4__21_), .B(regBoiz_regfile_5__21_), .S(
        net369145), .Z(n8454) );
  MUX2_X2 U12152 ( .A(regBoiz_regfile_6__21_), .B(regBoiz_regfile_7__21_), .S(
        net369147), .Z(n8453) );
  MUX2_X2 U12153 ( .A(n8454), .B(n8453), .S(n6804), .Z(n8455) );
  MUX2_X2 U12154 ( .A(n8456), .B(n8455), .S(n6825), .Z(n8464) );
  MUX2_X2 U12155 ( .A(regBoiz_regfile_8__21_), .B(regBoiz_regfile_9__21_), .S(
        net369244), .Z(n8458) );
  MUX2_X2 U12156 ( .A(regBoiz_regfile_10__21_), .B(regBoiz_regfile_11__21_), 
        .S(net369145), .Z(n8457) );
  MUX2_X2 U12157 ( .A(n8458), .B(n8457), .S(n6804), .Z(n8462) );
  MUX2_X2 U12158 ( .A(regBoiz_regfile_12__21_), .B(regBoiz_regfile_13__21_), 
        .S(net369228), .Z(n8460) );
  MUX2_X2 U12159 ( .A(regBoiz_regfile_14__21_), .B(regBoiz_regfile_15__21_), 
        .S(net369144), .Z(n8459) );
  MUX2_X2 U12160 ( .A(n8460), .B(n8459), .S(n6802), .Z(n8461) );
  MUX2_X2 U12161 ( .A(n8462), .B(n8461), .S(n6825), .Z(n8463) );
  MUX2_X2 U12162 ( .A(n8464), .B(n8463), .S(n6831), .Z(n8480) );
  MUX2_X2 U12163 ( .A(regBoiz_regfile_16__21_), .B(regBoiz_regfile_17__21_), 
        .S(net369161), .Z(n8466) );
  MUX2_X2 U12164 ( .A(regBoiz_regfile_18__21_), .B(regBoiz_regfile_19__21_), 
        .S(net369228), .Z(n8465) );
  MUX2_X2 U12165 ( .A(n8466), .B(n8465), .S(n6804), .Z(n8470) );
  MUX2_X2 U12166 ( .A(regBoiz_regfile_20__21_), .B(regBoiz_regfile_21__21_), 
        .S(net369145), .Z(n8468) );
  MUX2_X2 U12167 ( .A(regBoiz_regfile_22__21_), .B(regBoiz_regfile_23__21_), 
        .S(net369144), .Z(n8467) );
  MUX2_X2 U12168 ( .A(n8468), .B(n8467), .S(n6802), .Z(n8469) );
  MUX2_X2 U12169 ( .A(n8470), .B(n8469), .S(n6825), .Z(n8478) );
  MUX2_X2 U12170 ( .A(regBoiz_regfile_24__21_), .B(regBoiz_regfile_25__21_), 
        .S(net369162), .Z(n8472) );
  MUX2_X2 U12171 ( .A(regBoiz_regfile_26__21_), .B(regBoiz_regfile_27__21_), 
        .S(net369145), .Z(n8471) );
  MUX2_X2 U12172 ( .A(n8472), .B(n8471), .S(n6801), .Z(n8476) );
  MUX2_X2 U12173 ( .A(regBoiz_regfile_28__21_), .B(regBoiz_regfile_29__21_), 
        .S(net369220), .Z(n8474) );
  MUX2_X2 U12174 ( .A(regBoiz_regfile_30__21_), .B(regBoiz_regfile_31__21_), 
        .S(net377338), .Z(n8473) );
  MUX2_X2 U12175 ( .A(n8474), .B(n8473), .S(n6800), .Z(n8475) );
  MUX2_X2 U12176 ( .A(n8476), .B(n8475), .S(n6825), .Z(n8477) );
  MUX2_X2 U12177 ( .A(n8478), .B(n8477), .S(n6831), .Z(n8479) );
  MUX2_X2 U12178 ( .A(n8480), .B(n8479), .S(n6835), .Z(n12954) );
  NAND2_X2 U12179 ( .A1(n9718), .A2(n12954), .ZN(n8482) );
  NAND2_X2 U12180 ( .A1(daddr[10]), .A2(n6547), .ZN(n8481) );
  INV_X4 U12181 ( .A(n10417), .ZN(n9615) );
  XNOR2_X2 U12182 ( .A(n6565), .B(n9615), .ZN(n8484) );
  INV_X4 U12183 ( .A(n8484), .ZN(n8626) );
  NAND2_X2 U12184 ( .A1(n8626), .A2(net368519), .ZN(n9064) );
  NAND2_X2 U12185 ( .A1(aluBoi_imm32w_11_), .A2(n6556), .ZN(n8517) );
  MUX2_X2 U12186 ( .A(regBoiz_regfile_0__20_), .B(regBoiz_regfile_1__20_), .S(
        net378318), .Z(n8486) );
  MUX2_X2 U12187 ( .A(regBoiz_regfile_2__20_), .B(regBoiz_regfile_3__20_), .S(
        net377337), .Z(n8485) );
  MUX2_X2 U12188 ( .A(n8486), .B(n8485), .S(n6809), .Z(n8490) );
  MUX2_X2 U12189 ( .A(regBoiz_regfile_4__20_), .B(regBoiz_regfile_5__20_), .S(
        net369234), .Z(n8488) );
  MUX2_X2 U12190 ( .A(regBoiz_regfile_6__20_), .B(regBoiz_regfile_7__20_), .S(
        net369157), .Z(n8487) );
  MUX2_X2 U12191 ( .A(n8488), .B(n8487), .S(n6809), .Z(n8489) );
  MUX2_X2 U12192 ( .A(n8490), .B(n8489), .S(n6825), .Z(n8498) );
  MUX2_X2 U12193 ( .A(regBoiz_regfile_8__20_), .B(regBoiz_regfile_9__20_), .S(
        net369242), .Z(n8492) );
  MUX2_X2 U12194 ( .A(regBoiz_regfile_10__20_), .B(regBoiz_regfile_11__20_), 
        .S(net369166), .Z(n8491) );
  MUX2_X2 U12195 ( .A(n8492), .B(n8491), .S(n6809), .Z(n8496) );
  MUX2_X2 U12196 ( .A(regBoiz_regfile_12__20_), .B(regBoiz_regfile_13__20_), 
        .S(net369212), .Z(n8494) );
  MUX2_X2 U12197 ( .A(regBoiz_regfile_14__20_), .B(regBoiz_regfile_15__20_), 
        .S(net369226), .Z(n8493) );
  MUX2_X2 U12198 ( .A(n8494), .B(n8493), .S(n6809), .Z(n8495) );
  MUX2_X2 U12199 ( .A(n8496), .B(n8495), .S(n6825), .Z(n8497) );
  MUX2_X2 U12200 ( .A(n8498), .B(n8497), .S(n6831), .Z(n8514) );
  MUX2_X2 U12201 ( .A(regBoiz_regfile_16__20_), .B(regBoiz_regfile_17__20_), 
        .S(net369145), .Z(n8500) );
  MUX2_X2 U12202 ( .A(regBoiz_regfile_18__20_), .B(regBoiz_regfile_19__20_), 
        .S(net369220), .Z(n8499) );
  MUX2_X2 U12203 ( .A(n8500), .B(n8499), .S(n6809), .Z(n8504) );
  MUX2_X2 U12204 ( .A(regBoiz_regfile_20__20_), .B(regBoiz_regfile_21__20_), 
        .S(net369226), .Z(n8502) );
  MUX2_X2 U12205 ( .A(regBoiz_regfile_22__20_), .B(regBoiz_regfile_23__20_), 
        .S(net369163), .Z(n8501) );
  MUX2_X2 U12206 ( .A(n8502), .B(n8501), .S(n6809), .Z(n8503) );
  MUX2_X2 U12207 ( .A(n8504), .B(n8503), .S(n6825), .Z(n8512) );
  MUX2_X2 U12208 ( .A(regBoiz_regfile_24__20_), .B(regBoiz_regfile_25__20_), 
        .S(net369244), .Z(n8506) );
  MUX2_X2 U12209 ( .A(regBoiz_regfile_26__20_), .B(regBoiz_regfile_27__20_), 
        .S(net369166), .Z(n8505) );
  MUX2_X2 U12210 ( .A(n8506), .B(n8505), .S(n6809), .Z(n8510) );
  MUX2_X2 U12211 ( .A(regBoiz_regfile_28__20_), .B(regBoiz_regfile_29__20_), 
        .S(net369144), .Z(n8508) );
  MUX2_X2 U12212 ( .A(regBoiz_regfile_30__20_), .B(regBoiz_regfile_31__20_), 
        .S(net369236), .Z(n8507) );
  MUX2_X2 U12213 ( .A(n8508), .B(n8507), .S(n6809), .Z(n8509) );
  MUX2_X2 U12214 ( .A(n8510), .B(n8509), .S(n6825), .Z(n8511) );
  MUX2_X2 U12215 ( .A(n8512), .B(n8511), .S(n6831), .Z(n8513) );
  MUX2_X2 U12216 ( .A(n8514), .B(n8513), .S(n6835), .Z(n13079) );
  NAND2_X2 U12217 ( .A1(n9718), .A2(n13079), .ZN(n8516) );
  NAND2_X2 U12218 ( .A1(daddr[11]), .A2(n6547), .ZN(n8515) );
  INV_X4 U12219 ( .A(n10421), .ZN(n9651) );
  XNOR2_X2 U12220 ( .A(n6565), .B(n9651), .ZN(n8727) );
  INV_X4 U12221 ( .A(n8727), .ZN(n8518) );
  NAND2_X2 U12222 ( .A1(n8518), .A2(n6539), .ZN(n8726) );
  NAND2_X2 U12223 ( .A1(aluBoi_imm32w_8_), .A2(n6556), .ZN(n8551) );
  MUX2_X2 U12224 ( .A(regBoiz_regfile_0__23_), .B(regBoiz_regfile_1__23_), .S(
        net369242), .Z(n8520) );
  MUX2_X2 U12225 ( .A(regBoiz_regfile_2__23_), .B(regBoiz_regfile_3__23_), .S(
        net369226), .Z(n8519) );
  MUX2_X2 U12226 ( .A(n8520), .B(n8519), .S(n6809), .Z(n8524) );
  MUX2_X2 U12227 ( .A(regBoiz_regfile_4__23_), .B(regBoiz_regfile_5__23_), .S(
        net369234), .Z(n8522) );
  MUX2_X2 U12228 ( .A(regBoiz_regfile_6__23_), .B(regBoiz_regfile_7__23_), .S(
        net369155), .Z(n8521) );
  MUX2_X2 U12229 ( .A(n8522), .B(n8521), .S(n6809), .Z(n8523) );
  MUX2_X2 U12230 ( .A(n8524), .B(n8523), .S(n6825), .Z(n8532) );
  MUX2_X2 U12231 ( .A(regBoiz_regfile_8__23_), .B(regBoiz_regfile_9__23_), .S(
        net377338), .Z(n8526) );
  MUX2_X2 U12232 ( .A(regBoiz_regfile_10__23_), .B(regBoiz_regfile_11__23_), 
        .S(net369218), .Z(n8525) );
  MUX2_X2 U12233 ( .A(n8526), .B(n8525), .S(n6809), .Z(n8530) );
  MUX2_X2 U12234 ( .A(regBoiz_regfile_12__23_), .B(regBoiz_regfile_13__23_), 
        .S(net369154), .Z(n8528) );
  MUX2_X2 U12235 ( .A(n8528), .B(n8527), .S(n6810), .Z(n8529) );
  MUX2_X2 U12236 ( .A(n8530), .B(n8529), .S(n6825), .Z(n8531) );
  MUX2_X2 U12237 ( .A(n8532), .B(n8531), .S(n6831), .Z(n8548) );
  MUX2_X2 U12238 ( .A(regBoiz_regfile_16__23_), .B(regBoiz_regfile_17__23_), 
        .S(net369242), .Z(n8534) );
  MUX2_X2 U12239 ( .A(regBoiz_regfile_18__23_), .B(regBoiz_regfile_19__23_), 
        .S(net369147), .Z(n8533) );
  MUX2_X2 U12240 ( .A(n8534), .B(n8533), .S(n6810), .Z(n8538) );
  MUX2_X2 U12241 ( .A(regBoiz_regfile_20__23_), .B(regBoiz_regfile_21__23_), 
        .S(net369157), .Z(n8536) );
  MUX2_X2 U12242 ( .A(regBoiz_regfile_22__23_), .B(regBoiz_regfile_23__23_), 
        .S(net369157), .Z(n8535) );
  MUX2_X2 U12243 ( .A(n8536), .B(n8535), .S(n6810), .Z(n8537) );
  MUX2_X2 U12244 ( .A(n8538), .B(n8537), .S(n6825), .Z(n8546) );
  MUX2_X2 U12245 ( .A(regBoiz_regfile_24__23_), .B(regBoiz_regfile_25__23_), 
        .S(net369242), .Z(n8540) );
  MUX2_X2 U12246 ( .A(regBoiz_regfile_26__23_), .B(regBoiz_regfile_27__23_), 
        .S(net369214), .Z(n8539) );
  MUX2_X2 U12247 ( .A(n8540), .B(n8539), .S(n6810), .Z(n8544) );
  MUX2_X2 U12248 ( .A(regBoiz_regfile_28__23_), .B(regBoiz_regfile_29__23_), 
        .S(net369166), .Z(n8542) );
  MUX2_X2 U12249 ( .A(regBoiz_regfile_30__23_), .B(regBoiz_regfile_31__23_), 
        .S(net369144), .Z(n8541) );
  MUX2_X2 U12250 ( .A(n8542), .B(n8541), .S(n6810), .Z(n8543) );
  MUX2_X2 U12251 ( .A(n8544), .B(n8543), .S(n6825), .Z(n8545) );
  MUX2_X2 U12252 ( .A(n8546), .B(n8545), .S(n6831), .Z(n8547) );
  MUX2_X2 U12253 ( .A(n8548), .B(n8547), .S(n6835), .Z(n12988) );
  NAND2_X2 U12254 ( .A1(n9718), .A2(n12988), .ZN(n8550) );
  NAND2_X2 U12255 ( .A1(daddr[8]), .A2(n6547), .ZN(n8549) );
  INV_X4 U12256 ( .A(n10414), .ZN(n9625) );
  XNOR2_X2 U12257 ( .A(n6565), .B(n9625), .ZN(n8552) );
  INV_X4 U12258 ( .A(n8552), .ZN(n8588) );
  INV_X4 U12259 ( .A(n9075), .ZN(n8624) );
  NAND2_X2 U12260 ( .A1(aluBoi_imm32w_7_), .A2(n6556), .ZN(n8585) );
  MUX2_X2 U12261 ( .A(regBoiz_regfile_0__24_), .B(regBoiz_regfile_1__24_), .S(
        net369165), .Z(n8554) );
  MUX2_X2 U12262 ( .A(regBoiz_regfile_2__24_), .B(regBoiz_regfile_3__24_), .S(
        net369226), .Z(n8553) );
  MUX2_X2 U12263 ( .A(n8554), .B(n8553), .S(n6810), .Z(n8558) );
  MUX2_X2 U12264 ( .A(regBoiz_regfile_4__24_), .B(regBoiz_regfile_5__24_), .S(
        net369234), .Z(n8556) );
  MUX2_X2 U12265 ( .A(regBoiz_regfile_6__24_), .B(regBoiz_regfile_7__24_), .S(
        net369154), .Z(n8555) );
  MUX2_X2 U12266 ( .A(n8556), .B(n8555), .S(n6810), .Z(n8557) );
  MUX2_X2 U12267 ( .A(n8558), .B(n8557), .S(n6825), .Z(n8566) );
  MUX2_X2 U12268 ( .A(regBoiz_regfile_8__24_), .B(regBoiz_regfile_9__24_), .S(
        net377337), .Z(n8560) );
  MUX2_X2 U12269 ( .A(regBoiz_regfile_10__24_), .B(regBoiz_regfile_11__24_), 
        .S(net369246), .Z(n8559) );
  MUX2_X2 U12270 ( .A(n8560), .B(n8559), .S(n6810), .Z(n8564) );
  MUX2_X2 U12271 ( .A(regBoiz_regfile_12__24_), .B(regBoiz_regfile_13__24_), 
        .S(net369218), .Z(n8562) );
  MUX2_X2 U12272 ( .A(regBoiz_regfile_14__24_), .B(regBoiz_regfile_15__24_), 
        .S(net369165), .Z(n8561) );
  MUX2_X2 U12273 ( .A(n8562), .B(n8561), .S(n6810), .Z(n8563) );
  MUX2_X2 U12274 ( .A(n8564), .B(n8563), .S(n6825), .Z(n8565) );
  MUX2_X2 U12275 ( .A(n8566), .B(n8565), .S(n6831), .Z(n8582) );
  MUX2_X2 U12276 ( .A(regBoiz_regfile_16__24_), .B(regBoiz_regfile_17__24_), 
        .S(net369144), .Z(n8568) );
  MUX2_X2 U12277 ( .A(regBoiz_regfile_18__24_), .B(regBoiz_regfile_19__24_), 
        .S(net369165), .Z(n8567) );
  MUX2_X2 U12278 ( .A(n8568), .B(n8567), .S(n6810), .Z(n8572) );
  MUX2_X2 U12279 ( .A(regBoiz_regfile_20__24_), .B(regBoiz_regfile_21__24_), 
        .S(net369163), .Z(n8570) );
  MUX2_X2 U12280 ( .A(regBoiz_regfile_22__24_), .B(regBoiz_regfile_23__24_), 
        .S(net369214), .Z(n8569) );
  MUX2_X2 U12281 ( .A(n8570), .B(n8569), .S(n6810), .Z(n8571) );
  MUX2_X2 U12282 ( .A(n8572), .B(n8571), .S(n6824), .Z(n8580) );
  MUX2_X2 U12283 ( .A(regBoiz_regfile_24__24_), .B(regBoiz_regfile_25__24_), 
        .S(net369144), .Z(n8574) );
  MUX2_X2 U12284 ( .A(regBoiz_regfile_26__24_), .B(regBoiz_regfile_27__24_), 
        .S(net369163), .Z(n8573) );
  MUX2_X2 U12285 ( .A(n8574), .B(n8573), .S(n6810), .Z(n8578) );
  MUX2_X2 U12286 ( .A(regBoiz_regfile_28__24_), .B(regBoiz_regfile_29__24_), 
        .S(net369166), .Z(n8576) );
  MUX2_X2 U12287 ( .A(regBoiz_regfile_30__24_), .B(regBoiz_regfile_31__24_), 
        .S(net369226), .Z(n8575) );
  MUX2_X2 U12288 ( .A(n8576), .B(n8575), .S(n6811), .Z(n8577) );
  MUX2_X2 U12289 ( .A(n8578), .B(n8577), .S(n6824), .Z(n8579) );
  MUX2_X2 U12290 ( .A(n8580), .B(n8579), .S(n6831), .Z(n8581) );
  MUX2_X2 U12291 ( .A(n8582), .B(n8581), .S(n6835), .Z(n13025) );
  NAND2_X2 U12292 ( .A1(n9718), .A2(n13025), .ZN(n8584) );
  NAND2_X2 U12293 ( .A1(daddr[7]), .A2(n6547), .ZN(n8583) );
  INV_X4 U12294 ( .A(n9072), .ZN(n9104) );
  INV_X4 U12295 ( .A(n5007), .ZN(n10309) );
  XNOR2_X2 U12296 ( .A(n10309), .B(n8588), .ZN(n9103) );
  OAI21_X4 U12297 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9076) );
  INV_X4 U12298 ( .A(n13706), .ZN(n10850) );
  NAND2_X2 U12299 ( .A1(aluBoi_imm32w_9_), .A2(n6556), .ZN(n8621) );
  MUX2_X2 U12300 ( .A(regBoiz_regfile_0__22_), .B(regBoiz_regfile_1__22_), .S(
        net369244), .Z(n8590) );
  MUX2_X2 U12301 ( .A(regBoiz_regfile_2__22_), .B(regBoiz_regfile_3__22_), .S(
        net369165), .Z(n8589) );
  MUX2_X2 U12302 ( .A(n8590), .B(n8589), .S(n6811), .Z(n8594) );
  MUX2_X2 U12303 ( .A(regBoiz_regfile_4__22_), .B(regBoiz_regfile_5__22_), .S(
        net369156), .Z(n8592) );
  MUX2_X2 U12304 ( .A(regBoiz_regfile_6__22_), .B(regBoiz_regfile_7__22_), .S(
        net369164), .Z(n8591) );
  MUX2_X2 U12305 ( .A(n8592), .B(n8591), .S(n6811), .Z(n8593) );
  MUX2_X2 U12306 ( .A(n8594), .B(n8593), .S(n6824), .Z(n8602) );
  MUX2_X2 U12307 ( .A(regBoiz_regfile_8__22_), .B(regBoiz_regfile_9__22_), .S(
        net369157), .Z(n8596) );
  MUX2_X2 U12308 ( .A(n8596), .B(n8595), .S(n6811), .Z(n8600) );
  MUX2_X2 U12309 ( .A(regBoiz_regfile_12__22_), .B(regBoiz_regfile_13__22_), 
        .S(net369165), .Z(n8598) );
  MUX2_X2 U12310 ( .A(n8598), .B(n8597), .S(n6811), .Z(n8599) );
  MUX2_X2 U12311 ( .A(n8600), .B(n8599), .S(n6824), .Z(n8601) );
  MUX2_X2 U12312 ( .A(n8602), .B(n8601), .S(n6831), .Z(n8618) );
  MUX2_X2 U12313 ( .A(regBoiz_regfile_16__22_), .B(regBoiz_regfile_17__22_), 
        .S(net369155), .Z(n8604) );
  MUX2_X2 U12314 ( .A(regBoiz_regfile_18__22_), .B(regBoiz_regfile_19__22_), 
        .S(net369161), .Z(n8603) );
  MUX2_X2 U12315 ( .A(n8604), .B(n8603), .S(n6811), .Z(n8608) );
  MUX2_X2 U12316 ( .A(regBoiz_regfile_20__22_), .B(regBoiz_regfile_21__22_), 
        .S(net369165), .Z(n8606) );
  MUX2_X2 U12317 ( .A(regBoiz_regfile_22__22_), .B(regBoiz_regfile_23__22_), 
        .S(net369214), .Z(n8605) );
  MUX2_X2 U12318 ( .A(n8606), .B(n8605), .S(n6811), .Z(n8607) );
  MUX2_X2 U12319 ( .A(n8608), .B(n8607), .S(n6824), .Z(n8616) );
  MUX2_X2 U12320 ( .A(regBoiz_regfile_24__22_), .B(regBoiz_regfile_25__22_), 
        .S(net369163), .Z(n8610) );
  MUX2_X2 U12321 ( .A(regBoiz_regfile_26__22_), .B(regBoiz_regfile_27__22_), 
        .S(net369166), .Z(n8609) );
  MUX2_X2 U12322 ( .A(n8610), .B(n8609), .S(n6811), .Z(n8614) );
  MUX2_X2 U12323 ( .A(regBoiz_regfile_28__22_), .B(regBoiz_regfile_29__22_), 
        .S(net369165), .Z(n8612) );
  MUX2_X2 U12324 ( .A(regBoiz_regfile_30__22_), .B(regBoiz_regfile_31__22_), 
        .S(net369165), .Z(n8611) );
  MUX2_X2 U12325 ( .A(n8612), .B(n8611), .S(n6811), .Z(n8613) );
  MUX2_X2 U12326 ( .A(n8614), .B(n8613), .S(n6824), .Z(n8615) );
  MUX2_X2 U12327 ( .A(n8616), .B(n8615), .S(n6832), .Z(n8617) );
  MUX2_X2 U12328 ( .A(n8618), .B(n8617), .S(n6835), .Z(n12965) );
  NAND2_X2 U12329 ( .A1(n9718), .A2(n12965), .ZN(n8620) );
  NAND2_X2 U12330 ( .A1(daddr[9]), .A2(n6547), .ZN(n8619) );
  INV_X4 U12331 ( .A(n10413), .ZN(n9637) );
  XNOR2_X2 U12332 ( .A(n6565), .B(n9637), .ZN(n8622) );
  INV_X4 U12333 ( .A(n8622), .ZN(n8625) );
  XNOR2_X2 U12334 ( .A(n10850), .B(n8625), .ZN(n9078) );
  OAI21_X4 U12335 ( .B1(n8624), .B2(n8623), .A(n9078), .ZN(n9068) );
  NAND2_X2 U12336 ( .A1(n8625), .A2(n13706), .ZN(n9067) );
  INV_X4 U12337 ( .A(net368519), .ZN(net361808) );
  XNOR2_X2 U12338 ( .A(net361808), .B(n8626), .ZN(n9070) );
  INV_X4 U12339 ( .A(n9070), .ZN(n8627) );
  AOI21_X4 U12340 ( .B1(n9068), .B2(n9067), .A(n8627), .ZN(n8724) );
  NAND2_X2 U12341 ( .A1(n9075), .A2(n9067), .ZN(n8628) );
  NAND2_X2 U12342 ( .A1(aluBoi_imm32w_6_), .A2(n6556), .ZN(n8661) );
  MUX2_X2 U12343 ( .A(regBoiz_regfile_0__25_), .B(regBoiz_regfile_1__25_), .S(
        net369144), .Z(n8630) );
  MUX2_X2 U12344 ( .A(regBoiz_regfile_2__25_), .B(regBoiz_regfile_3__25_), .S(
        net369164), .Z(n8629) );
  MUX2_X2 U12345 ( .A(n8630), .B(n8629), .S(n6811), .Z(n8634) );
  MUX2_X2 U12346 ( .A(regBoiz_regfile_4__25_), .B(regBoiz_regfile_5__25_), .S(
        net369157), .Z(n8632) );
  MUX2_X2 U12347 ( .A(regBoiz_regfile_6__25_), .B(regBoiz_regfile_7__25_), .S(
        net369222), .Z(n8631) );
  MUX2_X2 U12348 ( .A(n8632), .B(n8631), .S(n6811), .Z(n8633) );
  MUX2_X2 U12349 ( .A(n8634), .B(n8633), .S(n6824), .Z(n8642) );
  MUX2_X2 U12350 ( .A(regBoiz_regfile_8__25_), .B(regBoiz_regfile_9__25_), .S(
        net369163), .Z(n8636) );
  MUX2_X2 U12351 ( .A(regBoiz_regfile_10__25_), .B(regBoiz_regfile_11__25_), 
        .S(net369144), .Z(n8635) );
  MUX2_X2 U12352 ( .A(n8636), .B(n8635), .S(n6811), .Z(n8640) );
  MUX2_X2 U12353 ( .A(regBoiz_regfile_12__25_), .B(regBoiz_regfile_13__25_), 
        .S(net369145), .Z(n8638) );
  MUX2_X2 U12354 ( .A(regBoiz_regfile_14__25_), .B(regBoiz_regfile_15__25_), 
        .S(net369218), .Z(n8637) );
  MUX2_X2 U12355 ( .A(n8638), .B(n8637), .S(n6812), .Z(n8639) );
  MUX2_X2 U12356 ( .A(n8640), .B(n8639), .S(n6824), .Z(n8641) );
  MUX2_X2 U12357 ( .A(n8642), .B(n8641), .S(n6832), .Z(n8658) );
  MUX2_X2 U12358 ( .A(regBoiz_regfile_16__25_), .B(regBoiz_regfile_17__25_), 
        .S(net369156), .Z(n8644) );
  MUX2_X2 U12359 ( .A(regBoiz_regfile_18__25_), .B(regBoiz_regfile_19__25_), 
        .S(net369164), .Z(n8643) );
  MUX2_X2 U12360 ( .A(n8644), .B(n8643), .S(n6812), .Z(n8648) );
  MUX2_X2 U12361 ( .A(regBoiz_regfile_20__25_), .B(regBoiz_regfile_21__25_), 
        .S(net369214), .Z(n8646) );
  MUX2_X2 U12362 ( .A(regBoiz_regfile_22__25_), .B(regBoiz_regfile_23__25_), 
        .S(net369145), .Z(n8645) );
  MUX2_X2 U12363 ( .A(n8646), .B(n8645), .S(n6812), .Z(n8647) );
  MUX2_X2 U12364 ( .A(n8648), .B(n8647), .S(n6824), .Z(n8656) );
  MUX2_X2 U12365 ( .A(regBoiz_regfile_24__25_), .B(regBoiz_regfile_25__25_), 
        .S(net369163), .Z(n8650) );
  MUX2_X2 U12366 ( .A(regBoiz_regfile_26__25_), .B(regBoiz_regfile_27__25_), 
        .S(net369144), .Z(n8649) );
  MUX2_X2 U12367 ( .A(n8650), .B(n8649), .S(n6812), .Z(n8654) );
  MUX2_X2 U12368 ( .A(regBoiz_regfile_28__25_), .B(regBoiz_regfile_29__25_), 
        .S(net369242), .Z(n8652) );
  MUX2_X2 U12369 ( .A(regBoiz_regfile_30__25_), .B(regBoiz_regfile_31__25_), 
        .S(net369145), .Z(n8651) );
  MUX2_X2 U12370 ( .A(n8652), .B(n8651), .S(n6812), .Z(n8653) );
  MUX2_X2 U12371 ( .A(n8654), .B(n8653), .S(n6824), .Z(n8655) );
  MUX2_X2 U12372 ( .A(n8656), .B(n8655), .S(n6832), .Z(n8657) );
  MUX2_X2 U12373 ( .A(n8658), .B(n8657), .S(n6835), .Z(n13036) );
  NAND2_X2 U12374 ( .A1(daddr[6]), .A2(n6547), .ZN(n8659) );
  XNOR2_X2 U12375 ( .A(n6565), .B(n9610), .ZN(n8696) );
  NAND2_X2 U12376 ( .A1(n8662), .A2(n6543), .ZN(n9102) );
  NAND2_X2 U12377 ( .A1(aluBoi_imm32w_5_), .A2(n6556), .ZN(n8695) );
  MUX2_X2 U12378 ( .A(regBoiz_regfile_0__26_), .B(regBoiz_regfile_1__26_), .S(
        net369156), .Z(n8664) );
  MUX2_X2 U12379 ( .A(regBoiz_regfile_2__26_), .B(regBoiz_regfile_3__26_), .S(
        net369161), .Z(n8663) );
  MUX2_X2 U12380 ( .A(n8664), .B(n8663), .S(n6812), .Z(n8668) );
  MUX2_X2 U12381 ( .A(regBoiz_regfile_4__26_), .B(regBoiz_regfile_5__26_), .S(
        net369214), .Z(n8666) );
  MUX2_X2 U12382 ( .A(regBoiz_regfile_6__26_), .B(regBoiz_regfile_7__26_), .S(
        net369166), .Z(n8665) );
  MUX2_X2 U12383 ( .A(n8666), .B(n8665), .S(n6812), .Z(n8667) );
  MUX2_X2 U12384 ( .A(n8668), .B(n8667), .S(n6824), .Z(n8676) );
  MUX2_X2 U12385 ( .A(regBoiz_regfile_8__26_), .B(regBoiz_regfile_9__26_), .S(
        net369157), .Z(n8670) );
  MUX2_X2 U12386 ( .A(regBoiz_regfile_10__26_), .B(regBoiz_regfile_11__26_), 
        .S(net369165), .Z(n8669) );
  MUX2_X2 U12387 ( .A(n8670), .B(n8669), .S(n6812), .Z(n8674) );
  MUX2_X2 U12388 ( .A(regBoiz_regfile_12__26_), .B(regBoiz_regfile_13__26_), 
        .S(net369165), .Z(n8672) );
  MUX2_X2 U12389 ( .A(regBoiz_regfile_14__26_), .B(regBoiz_regfile_15__26_), 
        .S(net369157), .Z(n8671) );
  MUX2_X2 U12390 ( .A(n8672), .B(n8671), .S(n6812), .Z(n8673) );
  MUX2_X2 U12391 ( .A(n8674), .B(n8673), .S(n6824), .Z(n8675) );
  MUX2_X2 U12392 ( .A(n8676), .B(n8675), .S(n6832), .Z(n8692) );
  MUX2_X2 U12393 ( .A(regBoiz_regfile_16__26_), .B(regBoiz_regfile_17__26_), 
        .S(net369154), .Z(n8678) );
  MUX2_X2 U12394 ( .A(regBoiz_regfile_18__26_), .B(regBoiz_regfile_19__26_), 
        .S(net369154), .Z(n8677) );
  MUX2_X2 U12395 ( .A(n8678), .B(n8677), .S(n6812), .Z(n8682) );
  MUX2_X2 U12396 ( .A(regBoiz_regfile_20__26_), .B(regBoiz_regfile_21__26_), 
        .S(net369218), .Z(n8680) );
  MUX2_X2 U12397 ( .A(regBoiz_regfile_22__26_), .B(regBoiz_regfile_23__26_), 
        .S(net369166), .Z(n8679) );
  MUX2_X2 U12398 ( .A(n8680), .B(n8679), .S(n6812), .Z(n8681) );
  MUX2_X2 U12399 ( .A(n8682), .B(n8681), .S(n6824), .Z(n8690) );
  MUX2_X2 U12400 ( .A(regBoiz_regfile_24__26_), .B(regBoiz_regfile_25__26_), 
        .S(net369155), .Z(n8684) );
  MUX2_X2 U12401 ( .A(regBoiz_regfile_26__26_), .B(regBoiz_regfile_27__26_), 
        .S(net369214), .Z(n8683) );
  MUX2_X2 U12402 ( .A(n8684), .B(n8683), .S(n6812), .Z(n8688) );
  MUX2_X2 U12403 ( .A(regBoiz_regfile_28__26_), .B(regBoiz_regfile_29__26_), 
        .S(net369157), .Z(n8686) );
  MUX2_X2 U12404 ( .A(n8686), .B(n8685), .S(n6813), .Z(n8687) );
  MUX2_X2 U12405 ( .A(n8688), .B(n8687), .S(n6824), .Z(n8689) );
  MUX2_X2 U12406 ( .A(n8690), .B(n8689), .S(n6832), .Z(n8691) );
  MUX2_X2 U12407 ( .A(n8692), .B(n8691), .S(n6835), .Z(n12969) );
  NAND2_X2 U12408 ( .A1(n9718), .A2(n12969), .ZN(n8694) );
  NAND2_X2 U12409 ( .A1(daddr[5]), .A2(n6547), .ZN(n8693) );
  XNOR2_X2 U12410 ( .A(n6565), .B(n9492), .ZN(n8719) );
  XNOR2_X2 U12411 ( .A(n8696), .B(n6543), .ZN(n9097) );
  XNOR2_X2 U12412 ( .A(n6565), .B(net362485), .ZN(n8703) );
  XNOR2_X2 U12413 ( .A(n8703), .B(n6618), .ZN(n9083) );
  OAI21_X4 U12414 ( .B1(n5954), .B2(n8882), .A(n9083), .ZN(n9089) );
  XNOR2_X2 U12415 ( .A(n6565), .B(n6618), .ZN(n8704) );
  NAND2_X2 U12416 ( .A1(n8704), .A2(net377611), .ZN(n9088) );
  INV_X4 U12417 ( .A(net368498), .ZN(net364246) );
  XNOR2_X2 U12418 ( .A(n8707), .B(n9677), .ZN(n8715) );
  XNOR2_X2 U12419 ( .A(n8712), .B(n8711), .ZN(n9678) );
  XNOR2_X2 U12420 ( .A(n8715), .B(net368498), .ZN(n9086) );
  OAI21_X4 U12421 ( .B1(net364246), .B2(n6072), .A(n8714), .ZN(n8876) );
  XNOR2_X2 U12422 ( .A(n6614), .B(n9677), .ZN(n8716) );
  XNOR2_X2 U12423 ( .A(n8716), .B(net368502), .ZN(n8875) );
  INV_X4 U12424 ( .A(n9088), .ZN(n8717) );
  NOR2_X4 U12425 ( .A1(n8717), .A2(n9087), .ZN(n8721) );
  NAND2_X2 U12426 ( .A1(n5021), .A2(n6545), .ZN(n8720) );
  OAI21_X4 U12427 ( .B1(n8721), .B2(n9093), .A(n8720), .ZN(n9094) );
  NAND4_X2 U12428 ( .A1(n9100), .A2(n9101), .A3(n8722), .A4(n9102), .ZN(n8723)
         );
  INV_X4 U12429 ( .A(n8725), .ZN(n8765) );
  INV_X4 U12430 ( .A(n8726), .ZN(n9464) );
  XNOR2_X2 U12431 ( .A(n8727), .B(n6539), .ZN(n9465) );
  NAND2_X2 U12432 ( .A1(aluBoi_imm32w_12_), .A2(n6556), .ZN(n8760) );
  MUX2_X2 U12433 ( .A(regBoiz_regfile_0__19_), .B(regBoiz_regfile_1__19_), .S(
        net369164), .Z(n8729) );
  MUX2_X2 U12434 ( .A(regBoiz_regfile_2__19_), .B(regBoiz_regfile_3__19_), .S(
        net369155), .Z(n8728) );
  MUX2_X2 U12435 ( .A(n8729), .B(n8728), .S(n6813), .Z(n8733) );
  MUX2_X2 U12436 ( .A(regBoiz_regfile_4__19_), .B(regBoiz_regfile_5__19_), .S(
        net369220), .Z(n8731) );
  MUX2_X2 U12437 ( .A(regBoiz_regfile_6__19_), .B(regBoiz_regfile_7__19_), .S(
        net369157), .Z(n8730) );
  MUX2_X2 U12438 ( .A(n8731), .B(n8730), .S(n6813), .Z(n8732) );
  MUX2_X2 U12439 ( .A(n8733), .B(n8732), .S(n6824), .Z(n8741) );
  MUX2_X2 U12440 ( .A(regBoiz_regfile_8__19_), .B(regBoiz_regfile_9__19_), .S(
        net369154), .Z(n8735) );
  MUX2_X2 U12441 ( .A(regBoiz_regfile_10__19_), .B(regBoiz_regfile_11__19_), 
        .S(net369228), .Z(n8734) );
  MUX2_X2 U12442 ( .A(n8735), .B(n8734), .S(n6813), .Z(n8739) );
  MUX2_X2 U12443 ( .A(regBoiz_regfile_12__19_), .B(regBoiz_regfile_13__19_), 
        .S(net369244), .Z(n8737) );
  MUX2_X2 U12444 ( .A(regBoiz_regfile_14__19_), .B(regBoiz_regfile_15__19_), 
        .S(net369244), .Z(n8736) );
  MUX2_X2 U12445 ( .A(n8737), .B(n8736), .S(n6813), .Z(n8738) );
  MUX2_X2 U12446 ( .A(n8739), .B(n8738), .S(n6824), .Z(n8740) );
  MUX2_X2 U12447 ( .A(n8741), .B(n8740), .S(n6831), .Z(n8757) );
  MUX2_X2 U12448 ( .A(regBoiz_regfile_16__19_), .B(regBoiz_regfile_17__19_), 
        .S(net369244), .Z(n8743) );
  MUX2_X2 U12449 ( .A(regBoiz_regfile_18__19_), .B(regBoiz_regfile_19__19_), 
        .S(net369234), .Z(n8742) );
  MUX2_X2 U12450 ( .A(n8743), .B(n8742), .S(n6813), .Z(n8747) );
  MUX2_X2 U12451 ( .A(regBoiz_regfile_20__19_), .B(regBoiz_regfile_21__19_), 
        .S(net369147), .Z(n8745) );
  MUX2_X2 U12452 ( .A(regBoiz_regfile_22__19_), .B(regBoiz_regfile_23__19_), 
        .S(net369242), .Z(n8744) );
  MUX2_X2 U12453 ( .A(n8745), .B(n8744), .S(n6813), .Z(n8746) );
  MUX2_X2 U12454 ( .A(n8747), .B(n8746), .S(n6824), .Z(n8755) );
  MUX2_X2 U12455 ( .A(regBoiz_regfile_24__19_), .B(regBoiz_regfile_25__19_), 
        .S(net377338), .Z(n8749) );
  MUX2_X2 U12456 ( .A(regBoiz_regfile_26__19_), .B(regBoiz_regfile_27__19_), 
        .S(net369234), .Z(n8748) );
  MUX2_X2 U12457 ( .A(n8749), .B(n8748), .S(n6813), .Z(n8753) );
  MUX2_X2 U12458 ( .A(regBoiz_regfile_28__19_), .B(regBoiz_regfile_29__19_), 
        .S(net369226), .Z(n8751) );
  MUX2_X2 U12459 ( .A(regBoiz_regfile_30__19_), .B(regBoiz_regfile_31__19_), 
        .S(net369156), .Z(n8750) );
  MUX2_X2 U12460 ( .A(n8751), .B(n8750), .S(n6813), .Z(n8752) );
  MUX2_X2 U12461 ( .A(n8753), .B(n8752), .S(n6824), .Z(n8754) );
  MUX2_X2 U12462 ( .A(n8755), .B(n8754), .S(n6832), .Z(n8756) );
  MUX2_X2 U12463 ( .A(n8757), .B(n8756), .S(n6835), .Z(n13067) );
  NAND2_X2 U12464 ( .A1(n9718), .A2(n13067), .ZN(n8759) );
  NAND2_X2 U12465 ( .A1(daddr[12]), .A2(n6547), .ZN(n8758) );
  INV_X4 U12466 ( .A(n10420), .ZN(n9664) );
  XNOR2_X2 U12467 ( .A(n6565), .B(n9664), .ZN(n8761) );
  INV_X4 U12468 ( .A(n8761), .ZN(n8762) );
  NAND2_X2 U12469 ( .A1(n8762), .A2(n6537), .ZN(n8763) );
  OAI21_X4 U12470 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n9469) );
  INV_X4 U12471 ( .A(n8766), .ZN(n9473) );
  INV_X4 U12472 ( .A(n8767), .ZN(n8768) );
  NAND2_X2 U12473 ( .A1(n6556), .A2(aluBoi_imm32w_15_), .ZN(n8801) );
  MUX2_X2 U12474 ( .A(regBoiz_regfile_0__16_), .B(regBoiz_regfile_1__16_), .S(
        net369147), .Z(n8770) );
  MUX2_X2 U12475 ( .A(regBoiz_regfile_2__16_), .B(regBoiz_regfile_3__16_), .S(
        net369220), .Z(n8769) );
  MUX2_X2 U12476 ( .A(n8770), .B(n8769), .S(n6813), .Z(n8774) );
  MUX2_X2 U12477 ( .A(regBoiz_regfile_4__16_), .B(regBoiz_regfile_5__16_), .S(
        net369228), .Z(n8772) );
  MUX2_X2 U12478 ( .A(regBoiz_regfile_6__16_), .B(regBoiz_regfile_7__16_), .S(
        net369147), .Z(n8771) );
  MUX2_X2 U12479 ( .A(n8772), .B(n8771), .S(n6813), .Z(n8773) );
  MUX2_X2 U12480 ( .A(n8774), .B(n8773), .S(n6824), .Z(n8782) );
  MUX2_X2 U12481 ( .A(regBoiz_regfile_8__16_), .B(regBoiz_regfile_9__16_), .S(
        net369244), .Z(n8776) );
  MUX2_X2 U12482 ( .A(regBoiz_regfile_10__16_), .B(regBoiz_regfile_11__16_), 
        .S(net369165), .Z(n8775) );
  MUX2_X2 U12483 ( .A(n8776), .B(n8775), .S(n6813), .Z(n8780) );
  MUX2_X2 U12484 ( .A(regBoiz_regfile_12__16_), .B(regBoiz_regfile_13__16_), 
        .S(net369163), .Z(n8778) );
  MUX2_X2 U12485 ( .A(regBoiz_regfile_14__16_), .B(regBoiz_regfile_15__16_), 
        .S(net369244), .Z(n8777) );
  MUX2_X2 U12486 ( .A(n8778), .B(n8777), .S(n6805), .Z(n8779) );
  MUX2_X2 U12487 ( .A(n8780), .B(n8779), .S(n6824), .Z(n8781) );
  MUX2_X2 U12488 ( .A(n8782), .B(n8781), .S(n6832), .Z(n8798) );
  MUX2_X2 U12489 ( .A(regBoiz_regfile_16__16_), .B(regBoiz_regfile_17__16_), 
        .S(net378318), .Z(n8784) );
  MUX2_X2 U12490 ( .A(regBoiz_regfile_18__16_), .B(regBoiz_regfile_19__16_), 
        .S(net369155), .Z(n8783) );
  MUX2_X2 U12491 ( .A(n8784), .B(n8783), .S(n6805), .Z(n8788) );
  MUX2_X2 U12492 ( .A(regBoiz_regfile_20__16_), .B(regBoiz_regfile_21__16_), 
        .S(net369154), .Z(n8786) );
  MUX2_X2 U12493 ( .A(regBoiz_regfile_22__16_), .B(regBoiz_regfile_23__16_), 
        .S(net369145), .Z(n8785) );
  MUX2_X2 U12494 ( .A(n8786), .B(n8785), .S(n6802), .Z(n8787) );
  MUX2_X2 U12495 ( .A(n8788), .B(n8787), .S(n6824), .Z(n8796) );
  MUX2_X2 U12496 ( .A(regBoiz_regfile_24__16_), .B(regBoiz_regfile_25__16_), 
        .S(net369156), .Z(n8790) );
  MUX2_X2 U12497 ( .A(regBoiz_regfile_26__16_), .B(regBoiz_regfile_27__16_), 
        .S(net369230), .Z(n8789) );
  MUX2_X2 U12498 ( .A(n8790), .B(n8789), .S(n6803), .Z(n8794) );
  MUX2_X2 U12499 ( .A(regBoiz_regfile_28__16_), .B(regBoiz_regfile_29__16_), 
        .S(net369234), .Z(n8792) );
  MUX2_X2 U12500 ( .A(regBoiz_regfile_30__16_), .B(regBoiz_regfile_31__16_), 
        .S(net377337), .Z(n8791) );
  MUX2_X2 U12501 ( .A(n8792), .B(n8791), .S(n6806), .Z(n8793) );
  MUX2_X2 U12502 ( .A(n8794), .B(n8793), .S(n6824), .Z(n8795) );
  MUX2_X2 U12503 ( .A(n8796), .B(n8795), .S(n6832), .Z(n8797) );
  MUX2_X2 U12504 ( .A(n8798), .B(n8797), .S(n6835), .Z(n12935) );
  NAND2_X2 U12505 ( .A1(n9718), .A2(n12935), .ZN(n8800) );
  NAND2_X2 U12506 ( .A1(daddr[15]), .A2(n6547), .ZN(n8799) );
  INV_X4 U12507 ( .A(n10422), .ZN(n9193) );
  XNOR2_X2 U12508 ( .A(n6565), .B(n9193), .ZN(n8802) );
  XNOR2_X2 U12509 ( .A(n8802), .B(n13527), .ZN(n9461) );
  NAND2_X2 U12510 ( .A1(n9462), .A2(n9461), .ZN(n9055) );
  INV_X4 U12511 ( .A(n8802), .ZN(n8803) );
  NAND2_X2 U12512 ( .A1(n8803), .A2(n13527), .ZN(n8929) );
  NAND2_X2 U12513 ( .A1(n9055), .A2(n8929), .ZN(n8872) );
  MUX2_X2 U12514 ( .A(regBoiz_regfile_0__15_), .B(regBoiz_regfile_1__15_), .S(
        net369147), .Z(n8805) );
  MUX2_X2 U12515 ( .A(regBoiz_regfile_2__15_), .B(regBoiz_regfile_3__15_), .S(
        net369154), .Z(n8804) );
  MUX2_X2 U12516 ( .A(n8805), .B(n8804), .S(n6803), .Z(n8809) );
  MUX2_X2 U12517 ( .A(regBoiz_regfile_4__15_), .B(regBoiz_regfile_5__15_), .S(
        net369236), .Z(n8807) );
  MUX2_X2 U12518 ( .A(regBoiz_regfile_6__15_), .B(regBoiz_regfile_7__15_), .S(
        net369214), .Z(n8806) );
  MUX2_X2 U12519 ( .A(n8807), .B(n8806), .S(n6799), .Z(n8808) );
  MUX2_X2 U12520 ( .A(n8809), .B(n8808), .S(n6824), .Z(n8817) );
  MUX2_X2 U12521 ( .A(regBoiz_regfile_8__15_), .B(regBoiz_regfile_9__15_), .S(
        net369218), .Z(n8811) );
  MUX2_X2 U12522 ( .A(regBoiz_regfile_10__15_), .B(regBoiz_regfile_11__15_), 
        .S(net369156), .Z(n8810) );
  MUX2_X2 U12523 ( .A(n8811), .B(n8810), .S(n6799), .Z(n8815) );
  MUX2_X2 U12524 ( .A(regBoiz_regfile_12__15_), .B(regBoiz_regfile_13__15_), 
        .S(net369157), .Z(n8813) );
  MUX2_X2 U12525 ( .A(regBoiz_regfile_14__15_), .B(regBoiz_regfile_15__15_), 
        .S(net369157), .Z(n8812) );
  MUX2_X2 U12526 ( .A(n8813), .B(n8812), .S(n6799), .Z(n8814) );
  MUX2_X2 U12527 ( .A(n8815), .B(n8814), .S(n6824), .Z(n8816) );
  MUX2_X2 U12528 ( .A(n8817), .B(n8816), .S(n6832), .Z(n8833) );
  MUX2_X2 U12529 ( .A(regBoiz_regfile_16__15_), .B(regBoiz_regfile_17__15_), 
        .S(net369226), .Z(n8819) );
  MUX2_X2 U12530 ( .A(regBoiz_regfile_18__15_), .B(regBoiz_regfile_19__15_), 
        .S(net369154), .Z(n8818) );
  MUX2_X2 U12531 ( .A(n8819), .B(n8818), .S(n6799), .Z(n8823) );
  MUX2_X2 U12532 ( .A(regBoiz_regfile_20__15_), .B(regBoiz_regfile_21__15_), 
        .S(net369218), .Z(n8821) );
  MUX2_X2 U12533 ( .A(regBoiz_regfile_22__15_), .B(regBoiz_regfile_23__15_), 
        .S(net369218), .Z(n8820) );
  MUX2_X2 U12534 ( .A(n8821), .B(n8820), .S(n6799), .Z(n8822) );
  MUX2_X2 U12535 ( .A(n8823), .B(n8822), .S(n6824), .Z(n8831) );
  MUX2_X2 U12536 ( .A(regBoiz_regfile_24__15_), .B(regBoiz_regfile_25__15_), 
        .S(net369155), .Z(n8825) );
  MUX2_X2 U12537 ( .A(regBoiz_regfile_26__15_), .B(regBoiz_regfile_27__15_), 
        .S(net369154), .Z(n8824) );
  MUX2_X2 U12538 ( .A(n8825), .B(n8824), .S(n6799), .Z(n8829) );
  MUX2_X2 U12539 ( .A(regBoiz_regfile_28__15_), .B(regBoiz_regfile_29__15_), 
        .S(net369155), .Z(n8827) );
  MUX2_X2 U12540 ( .A(regBoiz_regfile_30__15_), .B(regBoiz_regfile_31__15_), 
        .S(net369157), .Z(n8826) );
  MUX2_X2 U12541 ( .A(n8827), .B(n8826), .S(n6799), .Z(n8828) );
  MUX2_X2 U12542 ( .A(n8829), .B(n8828), .S(n6824), .Z(n8830) );
  MUX2_X2 U12543 ( .A(n8831), .B(n8830), .S(n6832), .Z(n8832) );
  MUX2_X2 U12544 ( .A(n8833), .B(n8832), .S(n6835), .Z(n13118) );
  NAND2_X2 U12545 ( .A1(n9718), .A2(n13118), .ZN(n8836) );
  NAND2_X2 U12546 ( .A1(aluBoi_imm32w_15_), .A2(idOut_31_), .ZN(n10043) );
  NAND2_X2 U12547 ( .A1(daddr[16]), .A2(n6547), .ZN(n8835) );
  INV_X4 U12548 ( .A(n10426), .ZN(n9588) );
  XNOR2_X2 U12549 ( .A(n6565), .B(n9588), .ZN(n8870) );
  XNOR2_X2 U12550 ( .A(n8870), .B(n6529), .ZN(n8888) );
  XNOR2_X2 U12551 ( .A(n8872), .B(n8888), .ZN(n13122) );
  INV_X4 U12552 ( .A(n6527), .ZN(n10189) );
  MUX2_X2 U12553 ( .A(regBoiz_regfile_0__14_), .B(regBoiz_regfile_1__14_), .S(
        net369244), .Z(n8838) );
  MUX2_X2 U12554 ( .A(regBoiz_regfile_2__14_), .B(regBoiz_regfile_3__14_), .S(
        net369226), .Z(n8837) );
  MUX2_X2 U12555 ( .A(n8838), .B(n8837), .S(n6799), .Z(n8842) );
  MUX2_X2 U12556 ( .A(regBoiz_regfile_4__14_), .B(regBoiz_regfile_5__14_), .S(
        net369234), .Z(n8840) );
  MUX2_X2 U12557 ( .A(regBoiz_regfile_6__14_), .B(regBoiz_regfile_7__14_), .S(
        net377337), .Z(n8839) );
  MUX2_X2 U12558 ( .A(n8840), .B(n8839), .S(n6799), .Z(n8841) );
  MUX2_X2 U12559 ( .A(n8842), .B(n8841), .S(n6824), .Z(n8850) );
  MUX2_X2 U12560 ( .A(regBoiz_regfile_8__14_), .B(regBoiz_regfile_9__14_), .S(
        net377338), .Z(n8844) );
  MUX2_X2 U12561 ( .A(regBoiz_regfile_10__14_), .B(regBoiz_regfile_11__14_), 
        .S(net369242), .Z(n8843) );
  MUX2_X2 U12562 ( .A(n8844), .B(n8843), .S(n6799), .Z(n8848) );
  MUX2_X2 U12563 ( .A(regBoiz_regfile_12__14_), .B(regBoiz_regfile_13__14_), 
        .S(net369236), .Z(n8846) );
  MUX2_X2 U12564 ( .A(regBoiz_regfile_14__14_), .B(regBoiz_regfile_15__14_), 
        .S(net369236), .Z(n8845) );
  MUX2_X2 U12565 ( .A(n8846), .B(n8845), .S(n6800), .Z(n8847) );
  MUX2_X2 U12566 ( .A(n8848), .B(n8847), .S(n6824), .Z(n8849) );
  MUX2_X2 U12567 ( .A(n8850), .B(n8849), .S(n6832), .Z(n8866) );
  MUX2_X2 U12568 ( .A(regBoiz_regfile_16__14_), .B(regBoiz_regfile_17__14_), 
        .S(net369244), .Z(n8852) );
  MUX2_X2 U12569 ( .A(regBoiz_regfile_18__14_), .B(regBoiz_regfile_19__14_), 
        .S(net369226), .Z(n8851) );
  MUX2_X2 U12570 ( .A(n8852), .B(n8851), .S(n6800), .Z(n8856) );
  MUX2_X2 U12571 ( .A(regBoiz_regfile_20__14_), .B(regBoiz_regfile_21__14_), 
        .S(net377338), .Z(n8854) );
  MUX2_X2 U12572 ( .A(regBoiz_regfile_22__14_), .B(regBoiz_regfile_23__14_), 
        .S(net369234), .Z(n8853) );
  MUX2_X2 U12573 ( .A(n8854), .B(n8853), .S(n6800), .Z(n8855) );
  MUX2_X2 U12574 ( .A(n8856), .B(n8855), .S(n6824), .Z(n8864) );
  MUX2_X2 U12575 ( .A(regBoiz_regfile_24__14_), .B(regBoiz_regfile_25__14_), 
        .S(net369147), .Z(n8858) );
  MUX2_X2 U12576 ( .A(regBoiz_regfile_26__14_), .B(regBoiz_regfile_27__14_), 
        .S(net377337), .Z(n8857) );
  MUX2_X2 U12577 ( .A(n8858), .B(n8857), .S(n6800), .Z(n8862) );
  MUX2_X2 U12578 ( .A(regBoiz_regfile_28__14_), .B(regBoiz_regfile_29__14_), 
        .S(net369226), .Z(n8860) );
  MUX2_X2 U12579 ( .A(regBoiz_regfile_30__14_), .B(regBoiz_regfile_31__14_), 
        .S(net369246), .Z(n8859) );
  MUX2_X2 U12580 ( .A(n8860), .B(n8859), .S(n6800), .Z(n8861) );
  MUX2_X2 U12581 ( .A(n8862), .B(n8861), .S(n6824), .Z(n8863) );
  MUX2_X2 U12582 ( .A(n8864), .B(n8863), .S(n6832), .Z(n8865) );
  MUX2_X2 U12583 ( .A(n8866), .B(n8865), .S(n6835), .Z(n13107) );
  NAND2_X2 U12584 ( .A1(n9718), .A2(n13107), .ZN(n8868) );
  NAND2_X2 U12585 ( .A1(daddr[17]), .A2(n6547), .ZN(n8867) );
  INV_X4 U12586 ( .A(n10425), .ZN(n9600) );
  XNOR2_X2 U12587 ( .A(n6565), .B(n9600), .ZN(n8869) );
  INV_X4 U12588 ( .A(n8869), .ZN(n8886) );
  XNOR2_X2 U12589 ( .A(n10189), .B(n8886), .ZN(n8887) );
  INV_X4 U12590 ( .A(n8887), .ZN(n8874) );
  INV_X4 U12591 ( .A(n8870), .ZN(n8871) );
  NAND2_X2 U12592 ( .A1(n8871), .A2(n6529), .ZN(n8928) );
  INV_X4 U12593 ( .A(n8928), .ZN(n8889) );
  AOI21_X4 U12594 ( .B1(n8872), .B2(n8888), .A(n8889), .ZN(n8873) );
  XNOR2_X2 U12595 ( .A(n8874), .B(n8873), .ZN(n13111) );
  NAND2_X2 U12596 ( .A1(n13122), .A2(n13111), .ZN(n9048) );
  INV_X4 U12597 ( .A(n8876), .ZN(n8877) );
  XNOR2_X2 U12598 ( .A(n8878), .B(n8877), .ZN(n13260) );
  INV_X4 U12599 ( .A(n8881), .ZN(n9082) );
  XNOR2_X2 U12600 ( .A(n8882), .B(n9082), .ZN(n13247) );
  NAND2_X2 U12601 ( .A1(n13260), .A2(n13248), .ZN(n9047) );
  INV_X4 U12602 ( .A(n9461), .ZN(n8885) );
  NOR2_X4 U12603 ( .A1(n8885), .A2(n8884), .ZN(n8926) );
  NAND2_X2 U12604 ( .A1(n8886), .A2(n6527), .ZN(n9058) );
  INV_X4 U12605 ( .A(n9058), .ZN(n8924) );
  OAI21_X4 U12606 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n9059) );
  INV_X4 U12607 ( .A(n9059), .ZN(n8923) );
  INV_X4 U12608 ( .A(n6525), .ZN(n10177) );
  MUX2_X2 U12609 ( .A(regBoiz_regfile_0__13_), .B(regBoiz_regfile_1__13_), .S(
        net369162), .Z(n8891) );
  MUX2_X2 U12610 ( .A(regBoiz_regfile_2__13_), .B(regBoiz_regfile_3__13_), .S(
        net369144), .Z(n8890) );
  MUX2_X2 U12611 ( .A(n8891), .B(n8890), .S(n6800), .Z(n8895) );
  MUX2_X2 U12612 ( .A(regBoiz_regfile_4__13_), .B(regBoiz_regfile_5__13_), .S(
        net369161), .Z(n8893) );
  MUX2_X2 U12613 ( .A(regBoiz_regfile_6__13_), .B(regBoiz_regfile_7__13_), .S(
        net377337), .Z(n8892) );
  MUX2_X2 U12614 ( .A(n8893), .B(n8892), .S(n6800), .Z(n8894) );
  MUX2_X2 U12615 ( .A(n8895), .B(n8894), .S(n6824), .Z(n8903) );
  MUX2_X2 U12616 ( .A(regBoiz_regfile_8__13_), .B(regBoiz_regfile_9__13_), .S(
        net369165), .Z(n8897) );
  MUX2_X2 U12617 ( .A(regBoiz_regfile_10__13_), .B(regBoiz_regfile_11__13_), 
        .S(net369244), .Z(n8896) );
  MUX2_X2 U12618 ( .A(n8897), .B(n8896), .S(n6800), .Z(n8901) );
  MUX2_X2 U12619 ( .A(regBoiz_regfile_12__13_), .B(regBoiz_regfile_13__13_), 
        .S(net369234), .Z(n8899) );
  MUX2_X2 U12620 ( .A(regBoiz_regfile_14__13_), .B(regBoiz_regfile_15__13_), 
        .S(net369156), .Z(n8898) );
  MUX2_X2 U12621 ( .A(n8899), .B(n8898), .S(n6800), .Z(n8900) );
  MUX2_X2 U12622 ( .A(n8901), .B(n8900), .S(n6823), .Z(n8902) );
  MUX2_X2 U12623 ( .A(n8903), .B(n8902), .S(n6831), .Z(n8919) );
  MUX2_X2 U12624 ( .A(regBoiz_regfile_16__13_), .B(regBoiz_regfile_17__13_), 
        .S(net369164), .Z(n8905) );
  MUX2_X2 U12625 ( .A(regBoiz_regfile_18__13_), .B(regBoiz_regfile_19__13_), 
        .S(net369162), .Z(n8904) );
  MUX2_X2 U12626 ( .A(n8905), .B(n8904), .S(n6800), .Z(n8909) );
  MUX2_X2 U12627 ( .A(regBoiz_regfile_20__13_), .B(regBoiz_regfile_21__13_), 
        .S(net369165), .Z(n8907) );
  MUX2_X2 U12628 ( .A(regBoiz_regfile_22__13_), .B(regBoiz_regfile_23__13_), 
        .S(net369154), .Z(n8906) );
  MUX2_X2 U12629 ( .A(n8907), .B(n8906), .S(n6800), .Z(n8908) );
  MUX2_X2 U12630 ( .A(n8909), .B(n8908), .S(n6823), .Z(n8917) );
  MUX2_X2 U12631 ( .A(regBoiz_regfile_24__13_), .B(regBoiz_regfile_25__13_), 
        .S(net369147), .Z(n8911) );
  MUX2_X2 U12632 ( .A(regBoiz_regfile_26__13_), .B(regBoiz_regfile_27__13_), 
        .S(net369155), .Z(n8910) );
  MUX2_X2 U12633 ( .A(n8911), .B(n8910), .S(n6800), .Z(n8915) );
  MUX2_X2 U12634 ( .A(regBoiz_regfile_28__13_), .B(regBoiz_regfile_29__13_), 
        .S(net369218), .Z(n8913) );
  MUX2_X2 U12635 ( .A(regBoiz_regfile_30__13_), .B(regBoiz_regfile_31__13_), 
        .S(net369244), .Z(n8912) );
  MUX2_X2 U12636 ( .A(n8913), .B(n8912), .S(n6801), .Z(n8914) );
  MUX2_X2 U12637 ( .A(n8915), .B(n8914), .S(n6823), .Z(n8916) );
  MUX2_X2 U12638 ( .A(n8917), .B(n8916), .S(n6831), .Z(n8918) );
  MUX2_X2 U12639 ( .A(n8919), .B(n8918), .S(n6835), .Z(n13097) );
  NAND2_X2 U12640 ( .A1(n9718), .A2(n13097), .ZN(n8921) );
  NAND2_X2 U12641 ( .A1(daddr[18]), .A2(n6547), .ZN(n8920) );
  INV_X4 U12642 ( .A(n10424), .ZN(n9515) );
  XNOR2_X2 U12643 ( .A(n5762), .B(n9515), .ZN(n8922) );
  INV_X4 U12644 ( .A(n8922), .ZN(n8927) );
  XNOR2_X2 U12645 ( .A(n10177), .B(n8927), .ZN(n9061) );
  OAI21_X4 U12646 ( .B1(n8924), .B2(n8923), .A(n9061), .ZN(n8925) );
  INV_X4 U12647 ( .A(n8925), .ZN(n8934) );
  NAND2_X2 U12648 ( .A1(n8926), .A2(n8934), .ZN(n9051) );
  INV_X4 U12649 ( .A(n9051), .ZN(n8932) );
  NAND2_X2 U12650 ( .A1(n8927), .A2(n6525), .ZN(n8937) );
  NAND2_X2 U12651 ( .A1(n8929), .A2(n8928), .ZN(n9056) );
  OAI21_X4 U12652 ( .B1(n8924), .B2(n9056), .A(n8934), .ZN(n8936) );
  NOR3_X4 U12653 ( .A1(n8933), .A2(n8932), .A3(n8931), .ZN(n8975) );
  NAND2_X2 U12654 ( .A1(n9051), .A2(n9052), .ZN(n8971) );
  NAND2_X2 U12655 ( .A1(n8937), .A2(n8936), .ZN(n9049) );
  INV_X4 U12656 ( .A(n6523), .ZN(n11380) );
  MUX2_X2 U12657 ( .A(regBoiz_regfile_0__12_), .B(regBoiz_regfile_1__12_), .S(
        net369162), .Z(n8939) );
  MUX2_X2 U12658 ( .A(regBoiz_regfile_2__12_), .B(regBoiz_regfile_3__12_), .S(
        net369157), .Z(n8938) );
  MUX2_X2 U12659 ( .A(n8939), .B(n8938), .S(n6801), .Z(n8943) );
  MUX2_X2 U12660 ( .A(regBoiz_regfile_4__12_), .B(regBoiz_regfile_5__12_), .S(
        net369155), .Z(n8941) );
  MUX2_X2 U12661 ( .A(regBoiz_regfile_6__12_), .B(regBoiz_regfile_7__12_), .S(
        net369163), .Z(n8940) );
  MUX2_X2 U12662 ( .A(n8941), .B(n8940), .S(n6801), .Z(n8942) );
  MUX2_X2 U12663 ( .A(n8943), .B(n8942), .S(n6823), .Z(n8951) );
  MUX2_X2 U12664 ( .A(regBoiz_regfile_8__12_), .B(regBoiz_regfile_9__12_), .S(
        net369156), .Z(n8945) );
  MUX2_X2 U12665 ( .A(regBoiz_regfile_10__12_), .B(regBoiz_regfile_11__12_), 
        .S(net369162), .Z(n8944) );
  MUX2_X2 U12666 ( .A(n8945), .B(n8944), .S(n6801), .Z(n8949) );
  MUX2_X2 U12667 ( .A(regBoiz_regfile_12__12_), .B(regBoiz_regfile_13__12_), 
        .S(net369165), .Z(n8947) );
  MUX2_X2 U12668 ( .A(regBoiz_regfile_14__12_), .B(regBoiz_regfile_15__12_), 
        .S(net369145), .Z(n8946) );
  MUX2_X2 U12669 ( .A(n8947), .B(n8946), .S(n6801), .Z(n8948) );
  MUX2_X2 U12670 ( .A(n8949), .B(n8948), .S(n6823), .Z(n8950) );
  MUX2_X2 U12671 ( .A(n8951), .B(n8950), .S(n6831), .Z(n8967) );
  MUX2_X2 U12672 ( .A(regBoiz_regfile_16__12_), .B(regBoiz_regfile_17__12_), 
        .S(net369154), .Z(n8953) );
  MUX2_X2 U12673 ( .A(regBoiz_regfile_18__12_), .B(regBoiz_regfile_19__12_), 
        .S(net369157), .Z(n8952) );
  MUX2_X2 U12674 ( .A(n8953), .B(n8952), .S(n6801), .Z(n8957) );
  MUX2_X2 U12675 ( .A(regBoiz_regfile_20__12_), .B(regBoiz_regfile_21__12_), 
        .S(net369156), .Z(n8955) );
  MUX2_X2 U12676 ( .A(regBoiz_regfile_22__12_), .B(regBoiz_regfile_23__12_), 
        .S(net369165), .Z(n8954) );
  MUX2_X2 U12677 ( .A(n8955), .B(n8954), .S(n6801), .Z(n8956) );
  MUX2_X2 U12678 ( .A(n8957), .B(n8956), .S(n6823), .Z(n8965) );
  MUX2_X2 U12679 ( .A(regBoiz_regfile_24__12_), .B(regBoiz_regfile_25__12_), 
        .S(net369212), .Z(n8959) );
  MUX2_X2 U12680 ( .A(regBoiz_regfile_26__12_), .B(regBoiz_regfile_27__12_), 
        .S(net369161), .Z(n8958) );
  MUX2_X2 U12681 ( .A(n8959), .B(n8958), .S(n6801), .Z(n8963) );
  MUX2_X2 U12682 ( .A(regBoiz_regfile_28__12_), .B(regBoiz_regfile_29__12_), 
        .S(net369144), .Z(n8961) );
  MUX2_X2 U12683 ( .A(regBoiz_regfile_30__12_), .B(regBoiz_regfile_31__12_), 
        .S(net369220), .Z(n8960) );
  MUX2_X2 U12684 ( .A(n8961), .B(n8960), .S(n6801), .Z(n8962) );
  MUX2_X2 U12685 ( .A(n8963), .B(n8962), .S(n6823), .Z(n8964) );
  MUX2_X2 U12686 ( .A(n8965), .B(n8964), .S(n6831), .Z(n8966) );
  MUX2_X2 U12687 ( .A(n8967), .B(n8966), .S(n6835), .Z(n12931) );
  NAND2_X2 U12688 ( .A1(n9718), .A2(n12931), .ZN(n8969) );
  NAND2_X2 U12689 ( .A1(daddr[19]), .A2(n6547), .ZN(n8968) );
  INV_X4 U12690 ( .A(n10423), .ZN(n9503) );
  XNOR2_X2 U12691 ( .A(n5762), .B(n9503), .ZN(n8970) );
  INV_X4 U12692 ( .A(n8970), .ZN(n8972) );
  XNOR2_X2 U12693 ( .A(n11380), .B(n8972), .ZN(n9053) );
  NAND2_X2 U12694 ( .A1(n8972), .A2(n6523), .ZN(n8973) );
  OAI21_X4 U12695 ( .B1(n8975), .B2(n8974), .A(n8973), .ZN(n9044) );
  INV_X4 U12696 ( .A(n6521), .ZN(n11487) );
  MUX2_X2 U12697 ( .A(regBoiz_regfile_0__11_), .B(regBoiz_regfile_1__11_), .S(
        net369147), .Z(n8977) );
  MUX2_X2 U12698 ( .A(regBoiz_regfile_2__11_), .B(regBoiz_regfile_3__11_), .S(
        net369163), .Z(n8976) );
  MUX2_X2 U12699 ( .A(n8977), .B(n8976), .S(n6801), .Z(n8981) );
  MUX2_X2 U12700 ( .A(regBoiz_regfile_4__11_), .B(regBoiz_regfile_5__11_), .S(
        net369157), .Z(n8979) );
  MUX2_X2 U12701 ( .A(regBoiz_regfile_6__11_), .B(regBoiz_regfile_7__11_), .S(
        net369244), .Z(n8978) );
  MUX2_X2 U12702 ( .A(n8979), .B(n8978), .S(n6801), .Z(n8980) );
  MUX2_X2 U12703 ( .A(n8981), .B(n8980), .S(n6823), .Z(n8989) );
  MUX2_X2 U12704 ( .A(regBoiz_regfile_8__11_), .B(regBoiz_regfile_9__11_), .S(
        net369212), .Z(n8983) );
  MUX2_X2 U12705 ( .A(regBoiz_regfile_10__11_), .B(regBoiz_regfile_11__11_), 
        .S(net377337), .Z(n8982) );
  MUX2_X2 U12706 ( .A(n8983), .B(n8982), .S(n6801), .Z(n8987) );
  MUX2_X2 U12707 ( .A(regBoiz_regfile_12__11_), .B(regBoiz_regfile_13__11_), 
        .S(net369228), .Z(n8985) );
  MUX2_X2 U12708 ( .A(regBoiz_regfile_14__11_), .B(regBoiz_regfile_15__11_), 
        .S(net369145), .Z(n8984) );
  MUX2_X2 U12709 ( .A(n8985), .B(n8984), .S(n6802), .Z(n8986) );
  MUX2_X2 U12710 ( .A(n8987), .B(n8986), .S(n6823), .Z(n8988) );
  MUX2_X2 U12711 ( .A(n8989), .B(n8988), .S(n6831), .Z(n9005) );
  MUX2_X2 U12712 ( .A(regBoiz_regfile_16__11_), .B(regBoiz_regfile_17__11_), 
        .S(net369220), .Z(n8991) );
  MUX2_X2 U12713 ( .A(regBoiz_regfile_18__11_), .B(regBoiz_regfile_19__11_), 
        .S(net369244), .Z(n8990) );
  MUX2_X2 U12714 ( .A(n8991), .B(n8990), .S(n6802), .Z(n8995) );
  MUX2_X2 U12715 ( .A(regBoiz_regfile_20__11_), .B(regBoiz_regfile_21__11_), 
        .S(net369147), .Z(n8993) );
  MUX2_X2 U12716 ( .A(regBoiz_regfile_22__11_), .B(regBoiz_regfile_23__11_), 
        .S(net369161), .Z(n8992) );
  MUX2_X2 U12717 ( .A(n8993), .B(n8992), .S(n6802), .Z(n8994) );
  MUX2_X2 U12718 ( .A(n8995), .B(n8994), .S(n6823), .Z(n9003) );
  MUX2_X2 U12719 ( .A(regBoiz_regfile_24__11_), .B(regBoiz_regfile_25__11_), 
        .S(net369236), .Z(n8997) );
  MUX2_X2 U12720 ( .A(regBoiz_regfile_26__11_), .B(regBoiz_regfile_27__11_), 
        .S(net369165), .Z(n8996) );
  MUX2_X2 U12721 ( .A(n8997), .B(n8996), .S(n6802), .Z(n9001) );
  MUX2_X2 U12722 ( .A(regBoiz_regfile_28__11_), .B(regBoiz_regfile_29__11_), 
        .S(net369144), .Z(n8999) );
  MUX2_X2 U12723 ( .A(regBoiz_regfile_30__11_), .B(regBoiz_regfile_31__11_), 
        .S(net369166), .Z(n8998) );
  MUX2_X2 U12724 ( .A(n8999), .B(n8998), .S(n6802), .Z(n9000) );
  MUX2_X2 U12725 ( .A(n9001), .B(n9000), .S(n6823), .Z(n9002) );
  MUX2_X2 U12726 ( .A(n9003), .B(n9002), .S(n6832), .Z(n9004) );
  MUX2_X2 U12727 ( .A(n9005), .B(n9004), .S(n6835), .Z(n12924) );
  NAND2_X2 U12728 ( .A1(n9718), .A2(n12924), .ZN(n9007) );
  NAND2_X2 U12729 ( .A1(daddr[20]), .A2(n6547), .ZN(n9006) );
  INV_X4 U12730 ( .A(n10427), .ZN(n9497) );
  XNOR2_X2 U12731 ( .A(n5762), .B(n9497), .ZN(n9008) );
  INV_X4 U12732 ( .A(n9008), .ZN(n9009) );
  XNOR2_X2 U12733 ( .A(n11487), .B(n9009), .ZN(n9045) );
  MUX2_X2 U12734 ( .A(regBoiz_regfile_0__10_), .B(regBoiz_regfile_1__10_), .S(
        net369212), .Z(n9011) );
  MUX2_X2 U12735 ( .A(regBoiz_regfile_2__10_), .B(regBoiz_regfile_3__10_), .S(
        net369228), .Z(n9010) );
  MUX2_X2 U12736 ( .A(n9011), .B(n9010), .S(n6802), .Z(n9015) );
  MUX2_X2 U12737 ( .A(regBoiz_regfile_4__10_), .B(regBoiz_regfile_5__10_), .S(
        net369236), .Z(n9013) );
  MUX2_X2 U12738 ( .A(regBoiz_regfile_6__10_), .B(regBoiz_regfile_7__10_), .S(
        net378318), .Z(n9012) );
  MUX2_X2 U12739 ( .A(n9013), .B(n9012), .S(n6802), .Z(n9014) );
  MUX2_X2 U12740 ( .A(n9015), .B(n9014), .S(n6823), .Z(n9023) );
  MUX2_X2 U12741 ( .A(regBoiz_regfile_8__10_), .B(regBoiz_regfile_9__10_), .S(
        net377338), .Z(n9017) );
  MUX2_X2 U12742 ( .A(regBoiz_regfile_10__10_), .B(regBoiz_regfile_11__10_), 
        .S(net369144), .Z(n9016) );
  MUX2_X2 U12743 ( .A(n9017), .B(n9016), .S(n6802), .Z(n9021) );
  MUX2_X2 U12744 ( .A(regBoiz_regfile_12__10_), .B(regBoiz_regfile_13__10_), 
        .S(net369145), .Z(n9019) );
  MUX2_X2 U12745 ( .A(n9019), .B(n9018), .S(n6802), .Z(n9020) );
  MUX2_X2 U12746 ( .A(n9021), .B(n9020), .S(n6823), .Z(n9022) );
  MUX2_X2 U12747 ( .A(n9023), .B(n9022), .S(n6831), .Z(n9039) );
  MUX2_X2 U12748 ( .A(regBoiz_regfile_16__10_), .B(regBoiz_regfile_17__10_), 
        .S(net369244), .Z(n9025) );
  MUX2_X2 U12749 ( .A(regBoiz_regfile_18__10_), .B(regBoiz_regfile_19__10_), 
        .S(net369164), .Z(n9024) );
  MUX2_X2 U12750 ( .A(n9025), .B(n9024), .S(n6802), .Z(n9029) );
  MUX2_X2 U12751 ( .A(regBoiz_regfile_20__10_), .B(regBoiz_regfile_21__10_), 
        .S(net369166), .Z(n9027) );
  MUX2_X2 U12752 ( .A(regBoiz_regfile_22__10_), .B(regBoiz_regfile_23__10_), 
        .S(net369154), .Z(n9026) );
  MUX2_X2 U12753 ( .A(n9027), .B(n9026), .S(n6802), .Z(n9028) );
  MUX2_X2 U12754 ( .A(n9029), .B(n9028), .S(n6823), .Z(n9037) );
  MUX2_X2 U12755 ( .A(regBoiz_regfile_24__10_), .B(regBoiz_regfile_25__10_), 
        .S(net369165), .Z(n9031) );
  MUX2_X2 U12756 ( .A(regBoiz_regfile_26__10_), .B(regBoiz_regfile_27__10_), 
        .S(net369155), .Z(n9030) );
  MUX2_X2 U12757 ( .A(n9031), .B(n9030), .S(n6802), .Z(n9035) );
  MUX2_X2 U12758 ( .A(regBoiz_regfile_28__10_), .B(regBoiz_regfile_29__10_), 
        .S(net369156), .Z(n9033) );
  MUX2_X2 U12759 ( .A(regBoiz_regfile_30__10_), .B(regBoiz_regfile_31__10_), 
        .S(net378318), .Z(n9032) );
  MUX2_X2 U12760 ( .A(n9033), .B(n9032), .S(n6803), .Z(n9034) );
  MUX2_X2 U12761 ( .A(n9035), .B(n9034), .S(n6823), .Z(n9036) );
  MUX2_X2 U12762 ( .A(n9037), .B(n9036), .S(n6831), .Z(n9038) );
  MUX2_X2 U12763 ( .A(n9039), .B(n9038), .S(n6834), .Z(n13136) );
  NAND2_X2 U12764 ( .A1(n9718), .A2(n13136), .ZN(n9041) );
  NAND2_X2 U12765 ( .A1(daddr[21]), .A2(n6547), .ZN(n9040) );
  INV_X4 U12766 ( .A(n10428), .ZN(n9486) );
  XNOR2_X2 U12767 ( .A(n5762), .B(n9486), .ZN(n9117) );
  INV_X4 U12768 ( .A(n9117), .ZN(n9042) );
  XNOR2_X2 U12769 ( .A(n11524), .B(n9042), .ZN(n9043) );
  INV_X4 U12770 ( .A(n9043), .ZN(n9115) );
  INV_X4 U12771 ( .A(n9049), .ZN(n9050) );
  OAI211_X2 U12772 ( .C1(n9473), .C2(n9052), .A(n9051), .B(n9050), .ZN(n9054)
         );
  XNOR2_X2 U12773 ( .A(n9054), .B(n9053), .ZN(n13090) );
  INV_X4 U12774 ( .A(n9055), .ZN(n9057) );
  NOR2_X4 U12775 ( .A1(n9057), .A2(n9056), .ZN(n9060) );
  OAI21_X4 U12776 ( .B1(n9060), .B2(n9059), .A(n9058), .ZN(n9062) );
  XNOR2_X2 U12777 ( .A(n9062), .B(n9061), .ZN(n13101) );
  INV_X4 U12778 ( .A(n13101), .ZN(n9063) );
  XNOR2_X2 U12779 ( .A(n9466), .B(n9465), .ZN(n13083) );
  XNOR2_X2 U12780 ( .A(n9071), .B(n9070), .ZN(n12958) );
  XNOR2_X2 U12781 ( .A(n9079), .B(n9078), .ZN(n12980) );
  XNOR2_X2 U12782 ( .A(n9084), .B(n9083), .ZN(n13010) );
  XNOR2_X2 U12783 ( .A(n9085), .B(n9086), .ZN(n13271) );
  XNOR2_X2 U12784 ( .A(n9099), .B(n9098), .ZN(n13040) );
  NAND4_X2 U12785 ( .A1(n13010), .A2(n13271), .A3(n12973), .A4(n13040), .ZN(
        n9110) );
  XNOR2_X2 U12786 ( .A(n9108), .B(n9107), .ZN(n13017) );
  NAND2_X2 U12787 ( .A1(n13029), .A2(n13017), .ZN(n9109) );
  MUX2_X2 U12788 ( .A(regBoiz_regfile_0__9_), .B(regBoiz_regfile_1__9_), .S(
        net369166), .Z(n9119) );
  MUX2_X2 U12789 ( .A(regBoiz_regfile_2__9_), .B(regBoiz_regfile_3__9_), .S(
        net377337), .Z(n9118) );
  MUX2_X2 U12790 ( .A(n9119), .B(n9118), .S(n6803), .Z(n9123) );
  MUX2_X2 U12791 ( .A(regBoiz_regfile_4__9_), .B(regBoiz_regfile_5__9_), .S(
        net369244), .Z(n9121) );
  MUX2_X2 U12792 ( .A(regBoiz_regfile_6__9_), .B(regBoiz_regfile_7__9_), .S(
        net369165), .Z(n9120) );
  MUX2_X2 U12793 ( .A(n9121), .B(n9120), .S(n6803), .Z(n9122) );
  MUX2_X2 U12794 ( .A(n9123), .B(n9122), .S(n6823), .Z(n9131) );
  MUX2_X2 U12795 ( .A(regBoiz_regfile_8__9_), .B(regBoiz_regfile_9__9_), .S(
        net369220), .Z(n9125) );
  MUX2_X2 U12796 ( .A(regBoiz_regfile_10__9_), .B(regBoiz_regfile_11__9_), .S(
        net369165), .Z(n9124) );
  MUX2_X2 U12797 ( .A(n9125), .B(n9124), .S(n6803), .Z(n9129) );
  MUX2_X2 U12798 ( .A(regBoiz_regfile_12__9_), .B(regBoiz_regfile_13__9_), .S(
        net369164), .Z(n9127) );
  MUX2_X2 U12799 ( .A(regBoiz_regfile_14__9_), .B(regBoiz_regfile_15__9_), .S(
        net369157), .Z(n9126) );
  MUX2_X2 U12800 ( .A(n9127), .B(n9126), .S(n6803), .Z(n9128) );
  MUX2_X2 U12801 ( .A(n9129), .B(n9128), .S(n6822), .Z(n9130) );
  MUX2_X2 U12802 ( .A(n9131), .B(n9130), .S(n6832), .Z(n9147) );
  MUX2_X2 U12803 ( .A(regBoiz_regfile_16__9_), .B(regBoiz_regfile_17__9_), .S(
        net369244), .Z(n9133) );
  MUX2_X2 U12804 ( .A(regBoiz_regfile_18__9_), .B(regBoiz_regfile_19__9_), .S(
        net369166), .Z(n9132) );
  MUX2_X2 U12805 ( .A(n9133), .B(n9132), .S(n6803), .Z(n9137) );
  MUX2_X2 U12806 ( .A(regBoiz_regfile_20__9_), .B(regBoiz_regfile_21__9_), .S(
        net369212), .Z(n9135) );
  MUX2_X2 U12807 ( .A(regBoiz_regfile_22__9_), .B(regBoiz_regfile_23__9_), .S(
        net369161), .Z(n9134) );
  MUX2_X2 U12808 ( .A(n9135), .B(n9134), .S(n6803), .Z(n9136) );
  MUX2_X2 U12809 ( .A(n9137), .B(n9136), .S(n6822), .Z(n9145) );
  MUX2_X2 U12810 ( .A(regBoiz_regfile_24__9_), .B(regBoiz_regfile_25__9_), .S(
        net369163), .Z(n9139) );
  MUX2_X2 U12811 ( .A(regBoiz_regfile_26__9_), .B(regBoiz_regfile_27__9_), .S(
        net369162), .Z(n9138) );
  MUX2_X2 U12812 ( .A(n9139), .B(n9138), .S(n6803), .Z(n9143) );
  MUX2_X2 U12813 ( .A(regBoiz_regfile_28__9_), .B(regBoiz_regfile_29__9_), .S(
        net369156), .Z(n9141) );
  MUX2_X2 U12814 ( .A(regBoiz_regfile_30__9_), .B(regBoiz_regfile_31__9_), .S(
        net369244), .Z(n9140) );
  MUX2_X2 U12815 ( .A(n9141), .B(n9140), .S(n6803), .Z(n9142) );
  MUX2_X2 U12816 ( .A(n9143), .B(n9142), .S(n6822), .Z(n9144) );
  MUX2_X2 U12817 ( .A(n9145), .B(n9144), .S(n6831), .Z(n9146) );
  MUX2_X2 U12818 ( .A(n9147), .B(n9146), .S(n6834), .Z(n13147) );
  NAND2_X2 U12819 ( .A1(n9718), .A2(n13147), .ZN(n9149) );
  NAND2_X2 U12820 ( .A1(daddr[22]), .A2(n6547), .ZN(n9148) );
  INV_X4 U12821 ( .A(n10429), .ZN(n9551) );
  XNOR2_X2 U12822 ( .A(n5762), .B(n9551), .ZN(n9150) );
  INV_X4 U12823 ( .A(n9150), .ZN(n9151) );
  XNOR2_X2 U12824 ( .A(net360723), .B(n9151), .ZN(n9200) );
  MUX2_X2 U12825 ( .A(regBoiz_regfile_0__8_), .B(regBoiz_regfile_1__8_), .S(
        net369244), .Z(n9153) );
  MUX2_X2 U12826 ( .A(regBoiz_regfile_2__8_), .B(regBoiz_regfile_3__8_), .S(
        net369164), .Z(n9152) );
  MUX2_X2 U12827 ( .A(n9153), .B(n9152), .S(n6803), .Z(n9157) );
  MUX2_X2 U12828 ( .A(regBoiz_regfile_4__8_), .B(regBoiz_regfile_5__8_), .S(
        net369165), .Z(n9155) );
  MUX2_X2 U12829 ( .A(regBoiz_regfile_6__8_), .B(regBoiz_regfile_7__8_), .S(
        net369212), .Z(n9154) );
  MUX2_X2 U12830 ( .A(n9155), .B(n9154), .S(n6803), .Z(n9156) );
  MUX2_X2 U12831 ( .A(n9157), .B(n9156), .S(n6822), .Z(n9165) );
  MUX2_X2 U12832 ( .A(regBoiz_regfile_8__8_), .B(regBoiz_regfile_9__8_), .S(
        net369163), .Z(n9159) );
  MUX2_X2 U12833 ( .A(regBoiz_regfile_10__8_), .B(regBoiz_regfile_11__8_), .S(
        net369161), .Z(n9158) );
  MUX2_X2 U12834 ( .A(n9159), .B(n9158), .S(n6803), .Z(n9163) );
  MUX2_X2 U12835 ( .A(regBoiz_regfile_12__8_), .B(regBoiz_regfile_13__8_), .S(
        net369156), .Z(n9161) );
  MUX2_X2 U12836 ( .A(regBoiz_regfile_14__8_), .B(regBoiz_regfile_15__8_), .S(
        net369228), .Z(n9160) );
  MUX2_X2 U12837 ( .A(n9161), .B(n9160), .S(n6804), .Z(n9162) );
  MUX2_X2 U12838 ( .A(n9163), .B(n9162), .S(n6822), .Z(n9164) );
  MUX2_X2 U12839 ( .A(n9165), .B(n9164), .S(n6831), .Z(n9181) );
  MUX2_X2 U12840 ( .A(regBoiz_regfile_16__8_), .B(regBoiz_regfile_17__8_), .S(
        net369157), .Z(n9167) );
  MUX2_X2 U12841 ( .A(regBoiz_regfile_18__8_), .B(regBoiz_regfile_19__8_), .S(
        net369155), .Z(n9166) );
  MUX2_X2 U12842 ( .A(n9167), .B(n9166), .S(n6804), .Z(n9171) );
  MUX2_X2 U12843 ( .A(regBoiz_regfile_20__8_), .B(regBoiz_regfile_21__8_), .S(
        net369154), .Z(n9169) );
  MUX2_X2 U12844 ( .A(regBoiz_regfile_22__8_), .B(regBoiz_regfile_23__8_), .S(
        net369236), .Z(n9168) );
  MUX2_X2 U12845 ( .A(n9169), .B(n9168), .S(n6804), .Z(n9170) );
  MUX2_X2 U12846 ( .A(n9171), .B(n9170), .S(n6822), .Z(n9179) );
  MUX2_X2 U12847 ( .A(regBoiz_regfile_24__8_), .B(regBoiz_regfile_25__8_), .S(
        net369156), .Z(n9173) );
  MUX2_X2 U12848 ( .A(regBoiz_regfile_26__8_), .B(regBoiz_regfile_27__8_), .S(
        net377338), .Z(n9172) );
  MUX2_X2 U12849 ( .A(n9173), .B(n9172), .S(n6804), .Z(n9177) );
  MUX2_X2 U12850 ( .A(regBoiz_regfile_28__8_), .B(regBoiz_regfile_29__8_), .S(
        net369228), .Z(n9175) );
  MUX2_X2 U12851 ( .A(regBoiz_regfile_30__8_), .B(regBoiz_regfile_31__8_), .S(
        net369165), .Z(n9174) );
  MUX2_X2 U12852 ( .A(n9175), .B(n9174), .S(n6804), .Z(n9176) );
  MUX2_X2 U12853 ( .A(n9177), .B(n9176), .S(n6822), .Z(n9178) );
  MUX2_X2 U12854 ( .A(n9179), .B(n9178), .S(n6831), .Z(n9180) );
  MUX2_X2 U12855 ( .A(n9181), .B(n9180), .S(n6834), .Z(n13157) );
  NAND2_X2 U12856 ( .A1(n9718), .A2(n13157), .ZN(n9183) );
  NAND2_X2 U12857 ( .A1(daddr[23]), .A2(n6547), .ZN(n9182) );
  INV_X4 U12858 ( .A(n10430), .ZN(n9565) );
  XNOR2_X2 U12859 ( .A(n5762), .B(n9565), .ZN(n9184) );
  INV_X4 U12860 ( .A(n9184), .ZN(n9377) );
  XNOR2_X2 U12861 ( .A(net360550), .B(n9377), .ZN(n9376) );
  NAND2_X2 U12862 ( .A1(aluBoi_aluBoi_shft_sraout[23]), .A2(n12944), .ZN(n9186) );
  NAND2_X2 U12863 ( .A1(aluBoi_aluBoi_shft_sllout[23]), .A2(n12940), .ZN(n9185) );
  INV_X4 U12864 ( .A(n13162), .ZN(n9206) );
  INV_X4 U12865 ( .A(n9188), .ZN(n9190) );
  NAND3_X4 U12866 ( .A1(n9190), .A2(n9189), .A3(n5345), .ZN(n9680) );
  MUX2_X2 U12867 ( .A(n9680), .B(n6564), .S(n9193), .Z(n9191) );
  NAND2_X2 U12868 ( .A1(n9191), .A2(n6561), .ZN(n9195) );
  INV_X4 U12869 ( .A(n13527), .ZN(n11316) );
  NAND2_X2 U12870 ( .A1(aluBoi_aluBoi_shft_srlout[15]), .A2(n6566), .ZN(n9197)
         );
  NAND2_X2 U12871 ( .A1(n9198), .A2(n9197), .ZN(n12946) );
  INV_X4 U12872 ( .A(n12946), .ZN(n9205) );
  NAND2_X2 U12873 ( .A1(aluBoi_aluBoi_shft_sraout[22]), .A2(n12944), .ZN(n9202) );
  NAND2_X2 U12874 ( .A1(aluBoi_aluBoi_shft_sllout[22]), .A2(n12940), .ZN(n9201) );
  NAND2_X2 U12875 ( .A1(aluBoi_aluBoi_shft_sllout[30]), .A2(n12940), .ZN(
        n13226) );
  NAND2_X2 U12876 ( .A1(aluBoi_aluBoi_shft_sraout[30]), .A2(n12944), .ZN(
        n13223) );
  NAND2_X2 U12877 ( .A1(n13226), .A2(n13223), .ZN(n9485) );
  MUX2_X2 U12878 ( .A(regBoiz_regfile_0__1_), .B(regBoiz_regfile_1__1_), .S(
        net369164), .Z(n9210) );
  MUX2_X2 U12879 ( .A(regBoiz_regfile_2__1_), .B(regBoiz_regfile_3__1_), .S(
        net369163), .Z(n9209) );
  MUX2_X2 U12880 ( .A(n9210), .B(n9209), .S(n6804), .Z(n9214) );
  MUX2_X2 U12881 ( .A(regBoiz_regfile_4__1_), .B(regBoiz_regfile_5__1_), .S(
        net369162), .Z(n9212) );
  MUX2_X2 U12882 ( .A(n9212), .B(n9211), .S(n6806), .Z(n9213) );
  MUX2_X2 U12883 ( .A(n9214), .B(n9213), .S(n6822), .Z(n9222) );
  MUX2_X2 U12884 ( .A(regBoiz_regfile_8__1_), .B(regBoiz_regfile_9__1_), .S(
        net369161), .Z(n9216) );
  MUX2_X2 U12885 ( .A(regBoiz_regfile_10__1_), .B(regBoiz_regfile_11__1_), .S(
        net369214), .Z(n9215) );
  MUX2_X2 U12886 ( .A(n9216), .B(n9215), .S(n6804), .Z(n9220) );
  MUX2_X2 U12887 ( .A(regBoiz_regfile_12__1_), .B(regBoiz_regfile_13__1_), .S(
        net369166), .Z(n9218) );
  MUX2_X2 U12888 ( .A(regBoiz_regfile_14__1_), .B(regBoiz_regfile_15__1_), .S(
        net369222), .Z(n9217) );
  MUX2_X2 U12889 ( .A(n9218), .B(n9217), .S(n6804), .Z(n9219) );
  MUX2_X2 U12890 ( .A(n9220), .B(n9219), .S(n6822), .Z(n9221) );
  MUX2_X2 U12891 ( .A(n9222), .B(n9221), .S(n6831), .Z(n9238) );
  MUX2_X2 U12892 ( .A(regBoiz_regfile_16__1_), .B(regBoiz_regfile_17__1_), .S(
        net369165), .Z(n9224) );
  MUX2_X2 U12893 ( .A(regBoiz_regfile_18__1_), .B(regBoiz_regfile_19__1_), .S(
        net369155), .Z(n9223) );
  MUX2_X2 U12894 ( .A(n9224), .B(n9223), .S(n6804), .Z(n9228) );
  MUX2_X2 U12895 ( .A(regBoiz_regfile_20__1_), .B(regBoiz_regfile_21__1_), .S(
        net369154), .Z(n9226) );
  MUX2_X2 U12896 ( .A(regBoiz_regfile_22__1_), .B(regBoiz_regfile_23__1_), .S(
        net377338), .Z(n9225) );
  MUX2_X2 U12897 ( .A(n9226), .B(n9225), .S(n6804), .Z(n9227) );
  MUX2_X2 U12898 ( .A(n9228), .B(n9227), .S(n6822), .Z(n9236) );
  MUX2_X2 U12899 ( .A(regBoiz_regfile_24__1_), .B(regBoiz_regfile_25__1_), .S(
        net369156), .Z(n9230) );
  MUX2_X2 U12900 ( .A(regBoiz_regfile_26__1_), .B(regBoiz_regfile_27__1_), .S(
        net369230), .Z(n9229) );
  MUX2_X2 U12901 ( .A(n9230), .B(n9229), .S(n6804), .Z(n9234) );
  MUX2_X2 U12902 ( .A(regBoiz_regfile_28__1_), .B(regBoiz_regfile_29__1_), .S(
        net369236), .Z(n9232) );
  MUX2_X2 U12903 ( .A(regBoiz_regfile_30__1_), .B(regBoiz_regfile_31__1_), .S(
        net377337), .Z(n9231) );
  MUX2_X2 U12904 ( .A(n9232), .B(n9231), .S(n6804), .Z(n9233) );
  MUX2_X2 U12905 ( .A(n9234), .B(n9233), .S(n6824), .Z(n9235) );
  MUX2_X2 U12906 ( .A(n9236), .B(n9235), .S(n6832), .Z(n9237) );
  MUX2_X2 U12907 ( .A(n9238), .B(n9237), .S(n6834), .Z(n13215) );
  NAND2_X2 U12908 ( .A1(n9718), .A2(n13215), .ZN(n9240) );
  NAND2_X2 U12909 ( .A1(daddr[30]), .A2(n6547), .ZN(n9239) );
  INV_X4 U12910 ( .A(n12312), .ZN(n9576) );
  XNOR2_X2 U12911 ( .A(n5762), .B(n9576), .ZN(n9728) );
  XNOR2_X2 U12912 ( .A(n9728), .B(n6509), .ZN(n13219) );
  MUX2_X2 U12913 ( .A(regBoiz_regfile_0__2_), .B(regBoiz_regfile_1__2_), .S(
        net378318), .Z(n9242) );
  MUX2_X2 U12914 ( .A(regBoiz_regfile_2__2_), .B(regBoiz_regfile_3__2_), .S(
        net369162), .Z(n9241) );
  MUX2_X2 U12915 ( .A(n9242), .B(n9241), .S(n6804), .Z(n9246) );
  MUX2_X2 U12916 ( .A(regBoiz_regfile_4__2_), .B(regBoiz_regfile_5__2_), .S(
        net369157), .Z(n9244) );
  MUX2_X2 U12917 ( .A(regBoiz_regfile_6__2_), .B(regBoiz_regfile_7__2_), .S(
        net369165), .Z(n9243) );
  MUX2_X2 U12918 ( .A(n9244), .B(n9243), .S(n6804), .Z(n9245) );
  MUX2_X2 U12919 ( .A(n9246), .B(n9245), .S(n6822), .Z(n9254) );
  MUX2_X2 U12920 ( .A(regBoiz_regfile_8__2_), .B(regBoiz_regfile_9__2_), .S(
        net369161), .Z(n9248) );
  MUX2_X2 U12921 ( .A(regBoiz_regfile_10__2_), .B(regBoiz_regfile_11__2_), .S(
        net369164), .Z(n9247) );
  MUX2_X2 U12922 ( .A(n9248), .B(n9247), .S(n6804), .Z(n9252) );
  MUX2_X2 U12923 ( .A(regBoiz_regfile_12__2_), .B(regBoiz_regfile_13__2_), .S(
        net369163), .Z(n9250) );
  MUX2_X2 U12924 ( .A(regBoiz_regfile_14__2_), .B(regBoiz_regfile_15__2_), .S(
        net369244), .Z(n9249) );
  MUX2_X2 U12925 ( .A(n9250), .B(n9249), .S(n6804), .Z(n9251) );
  MUX2_X2 U12926 ( .A(n9252), .B(n9251), .S(n6822), .Z(n9253) );
  MUX2_X2 U12927 ( .A(n9254), .B(n9253), .S(n6831), .Z(n9270) );
  MUX2_X2 U12928 ( .A(regBoiz_regfile_16__2_), .B(regBoiz_regfile_17__2_), .S(
        net369165), .Z(n9256) );
  MUX2_X2 U12929 ( .A(regBoiz_regfile_18__2_), .B(regBoiz_regfile_19__2_), .S(
        net369162), .Z(n9255) );
  MUX2_X2 U12930 ( .A(n9256), .B(n9255), .S(n6804), .Z(n9260) );
  MUX2_X2 U12931 ( .A(regBoiz_regfile_20__2_), .B(regBoiz_regfile_21__2_), .S(
        net369212), .Z(n9258) );
  MUX2_X2 U12932 ( .A(regBoiz_regfile_22__2_), .B(regBoiz_regfile_23__2_), .S(
        net369222), .Z(n9257) );
  MUX2_X2 U12933 ( .A(n9258), .B(n9257), .S(n6804), .Z(n9259) );
  MUX2_X2 U12934 ( .A(n9260), .B(n9259), .S(n6822), .Z(n9268) );
  MUX2_X2 U12935 ( .A(regBoiz_regfile_24__2_), .B(regBoiz_regfile_25__2_), .S(
        net369161), .Z(n9262) );
  MUX2_X2 U12936 ( .A(regBoiz_regfile_26__2_), .B(regBoiz_regfile_27__2_), .S(
        net377338), .Z(n9261) );
  MUX2_X2 U12937 ( .A(n9262), .B(n9261), .S(n6804), .Z(n9266) );
  MUX2_X2 U12938 ( .A(regBoiz_regfile_28__2_), .B(regBoiz_regfile_29__2_), .S(
        net369228), .Z(n9264) );
  MUX2_X2 U12939 ( .A(regBoiz_regfile_30__2_), .B(regBoiz_regfile_31__2_), .S(
        net369144), .Z(n9263) );
  MUX2_X2 U12940 ( .A(n9264), .B(n9263), .S(n6804), .Z(n9265) );
  MUX2_X2 U12941 ( .A(n9266), .B(n9265), .S(n6822), .Z(n9267) );
  MUX2_X2 U12942 ( .A(n9268), .B(n9267), .S(n6831), .Z(n9269) );
  MUX2_X2 U12943 ( .A(n9270), .B(n9269), .S(n6834), .Z(n13233) );
  NAND2_X2 U12944 ( .A1(n9718), .A2(n13233), .ZN(n9272) );
  NAND2_X2 U12945 ( .A1(daddr[29]), .A2(n6547), .ZN(n9271) );
  INV_X4 U12946 ( .A(n12491), .ZN(n9595) );
  XNOR2_X2 U12947 ( .A(n5762), .B(n9595), .ZN(n9456) );
  INV_X4 U12948 ( .A(n9456), .ZN(n9273) );
  XNOR2_X2 U12949 ( .A(n12249), .B(n9273), .ZN(n9743) );
  MUX2_X2 U12950 ( .A(regBoiz_regfile_0__3_), .B(regBoiz_regfile_1__3_), .S(
        net369220), .Z(n9275) );
  MUX2_X2 U12951 ( .A(regBoiz_regfile_2__3_), .B(regBoiz_regfile_3__3_), .S(
        net369244), .Z(n9274) );
  MUX2_X2 U12952 ( .A(n9275), .B(n9274), .S(n6804), .Z(n9279) );
  MUX2_X2 U12953 ( .A(regBoiz_regfile_4__3_), .B(regBoiz_regfile_5__3_), .S(
        net378318), .Z(n9277) );
  MUX2_X2 U12954 ( .A(regBoiz_regfile_6__3_), .B(regBoiz_regfile_7__3_), .S(
        net369164), .Z(n9276) );
  MUX2_X2 U12955 ( .A(n9277), .B(n9276), .S(n6804), .Z(n9278) );
  MUX2_X2 U12956 ( .A(n9279), .B(n9278), .S(n6822), .Z(n9287) );
  MUX2_X2 U12957 ( .A(regBoiz_regfile_8__3_), .B(regBoiz_regfile_9__3_), .S(
        net369147), .Z(n9281) );
  MUX2_X2 U12958 ( .A(regBoiz_regfile_10__3_), .B(regBoiz_regfile_11__3_), .S(
        net369212), .Z(n9280) );
  MUX2_X2 U12959 ( .A(n9281), .B(n9280), .S(n6804), .Z(n9285) );
  MUX2_X2 U12960 ( .A(regBoiz_regfile_12__3_), .B(regBoiz_regfile_13__3_), .S(
        net369165), .Z(n9283) );
  MUX2_X2 U12961 ( .A(regBoiz_regfile_14__3_), .B(regBoiz_regfile_15__3_), .S(
        net369154), .Z(n9282) );
  MUX2_X2 U12962 ( .A(n9283), .B(n9282), .S(n6804), .Z(n9284) );
  MUX2_X2 U12963 ( .A(n9285), .B(n9284), .S(n6822), .Z(n9286) );
  MUX2_X2 U12964 ( .A(n9287), .B(n9286), .S(n6831), .Z(n9303) );
  MUX2_X2 U12965 ( .A(regBoiz_regfile_16__3_), .B(regBoiz_regfile_17__3_), .S(
        net369145), .Z(n9289) );
  MUX2_X2 U12966 ( .A(regBoiz_regfile_18__3_), .B(regBoiz_regfile_19__3_), .S(
        net369155), .Z(n9288) );
  MUX2_X2 U12967 ( .A(n9289), .B(n9288), .S(n6804), .Z(n9293) );
  MUX2_X2 U12968 ( .A(regBoiz_regfile_20__3_), .B(regBoiz_regfile_21__3_), .S(
        net369154), .Z(n9291) );
  MUX2_X2 U12969 ( .A(regBoiz_regfile_22__3_), .B(regBoiz_regfile_23__3_), .S(
        net369230), .Z(n9290) );
  MUX2_X2 U12970 ( .A(n9291), .B(n9290), .S(n6804), .Z(n9292) );
  MUX2_X2 U12971 ( .A(n9293), .B(n9292), .S(n6823), .Z(n9301) );
  MUX2_X2 U12972 ( .A(regBoiz_regfile_24__3_), .B(regBoiz_regfile_25__3_), .S(
        net369156), .Z(n9295) );
  MUX2_X2 U12973 ( .A(regBoiz_regfile_26__3_), .B(regBoiz_regfile_27__3_), .S(
        net369236), .Z(n9294) );
  MUX2_X2 U12974 ( .A(n9295), .B(n9294), .S(n6804), .Z(n9299) );
  MUX2_X2 U12975 ( .A(regBoiz_regfile_28__3_), .B(regBoiz_regfile_29__3_), .S(
        net369220), .Z(n9297) );
  MUX2_X2 U12976 ( .A(regBoiz_regfile_30__3_), .B(regBoiz_regfile_31__3_), .S(
        net369165), .Z(n9296) );
  MUX2_X2 U12977 ( .A(n9297), .B(n9296), .S(n6804), .Z(n9298) );
  MUX2_X2 U12978 ( .A(n9299), .B(n9298), .S(n6823), .Z(n9300) );
  MUX2_X2 U12979 ( .A(n9301), .B(n9300), .S(n6832), .Z(n9302) );
  MUX2_X2 U12980 ( .A(n9303), .B(n9302), .S(n6835), .Z(n13187) );
  NAND2_X2 U12981 ( .A1(n9718), .A2(n13187), .ZN(n9305) );
  NAND2_X2 U12982 ( .A1(daddr[28]), .A2(n6547), .ZN(n9304) );
  INV_X4 U12983 ( .A(n12211), .ZN(n9530) );
  XNOR2_X2 U12984 ( .A(n5762), .B(n9530), .ZN(n9306) );
  XNOR2_X2 U12985 ( .A(n9306), .B(n6513), .ZN(n9761) );
  INV_X4 U12986 ( .A(n9761), .ZN(n9308) );
  INV_X4 U12987 ( .A(n9306), .ZN(n9307) );
  NAND2_X2 U12988 ( .A1(n9307), .A2(n6513), .ZN(n9742) );
  NAND2_X2 U12989 ( .A1(n9308), .A2(n9742), .ZN(n9455) );
  MUX2_X2 U12990 ( .A(regBoiz_regfile_0__4_), .B(regBoiz_regfile_1__4_), .S(
        net369144), .Z(n9310) );
  MUX2_X2 U12991 ( .A(regBoiz_regfile_2__4_), .B(regBoiz_regfile_3__4_), .S(
        net369166), .Z(n9309) );
  MUX2_X2 U12992 ( .A(n9310), .B(n9309), .S(n6804), .Z(n9314) );
  MUX2_X2 U12993 ( .A(regBoiz_regfile_4__4_), .B(regBoiz_regfile_5__4_), .S(
        net369155), .Z(n9312) );
  MUX2_X2 U12994 ( .A(n9312), .B(n9311), .S(n6804), .Z(n9313) );
  MUX2_X2 U12995 ( .A(n9314), .B(n9313), .S(n6822), .Z(n9322) );
  MUX2_X2 U12996 ( .A(regBoiz_regfile_8__4_), .B(regBoiz_regfile_9__4_), .S(
        net369156), .Z(n9316) );
  MUX2_X2 U12997 ( .A(n9316), .B(n9315), .S(n6804), .Z(n9320) );
  MUX2_X2 U12998 ( .A(regBoiz_regfile_12__4_), .B(regBoiz_regfile_13__4_), .S(
        net369236), .Z(n9318) );
  MUX2_X2 U12999 ( .A(n9318), .B(n9317), .S(n6804), .Z(n9319) );
  MUX2_X2 U13000 ( .A(n9320), .B(n9319), .S(n6823), .Z(n9321) );
  MUX2_X2 U13001 ( .A(n9322), .B(n9321), .S(n6832), .Z(n9338) );
  MUX2_X2 U13002 ( .A(regBoiz_regfile_16__4_), .B(regBoiz_regfile_17__4_), .S(
        net369154), .Z(n9324) );
  MUX2_X2 U13003 ( .A(regBoiz_regfile_18__4_), .B(regBoiz_regfile_19__4_), .S(
        net369145), .Z(n9323) );
  MUX2_X2 U13004 ( .A(n9324), .B(n9323), .S(n6804), .Z(n9328) );
  MUX2_X2 U13005 ( .A(regBoiz_regfile_20__4_), .B(regBoiz_regfile_21__4_), .S(
        net369236), .Z(n9326) );
  MUX2_X2 U13006 ( .A(regBoiz_regfile_22__4_), .B(regBoiz_regfile_23__4_), .S(
        net369163), .Z(n9325) );
  MUX2_X2 U13007 ( .A(n9326), .B(n9325), .S(n6804), .Z(n9327) );
  MUX2_X2 U13008 ( .A(n9328), .B(n9327), .S(n6825), .Z(n9336) );
  MUX2_X2 U13009 ( .A(regBoiz_regfile_24__4_), .B(regBoiz_regfile_25__4_), .S(
        net378318), .Z(n9330) );
  MUX2_X2 U13010 ( .A(n9330), .B(n9329), .S(n6804), .Z(n9334) );
  MUX2_X2 U13011 ( .A(regBoiz_regfile_28__4_), .B(regBoiz_regfile_29__4_), .S(
        net369157), .Z(n9332) );
  MUX2_X2 U13012 ( .A(regBoiz_regfile_30__4_), .B(regBoiz_regfile_31__4_), .S(
        net369147), .Z(n9331) );
  MUX2_X2 U13013 ( .A(n9332), .B(n9331), .S(n6805), .Z(n9333) );
  MUX2_X2 U13014 ( .A(n9334), .B(n9333), .S(n6823), .Z(n9335) );
  MUX2_X2 U13015 ( .A(n9336), .B(n9335), .S(n6830), .Z(n9337) );
  MUX2_X2 U13016 ( .A(n9338), .B(n9337), .S(n6834), .Z(n13195) );
  NAND2_X2 U13017 ( .A1(n9718), .A2(n13195), .ZN(n9340) );
  NAND2_X2 U13018 ( .A1(daddr[27]), .A2(n6547), .ZN(n9339) );
  INV_X4 U13019 ( .A(n10431), .ZN(n9545) );
  XNOR2_X2 U13020 ( .A(n5762), .B(n9545), .ZN(n9341) );
  INV_X4 U13021 ( .A(n9341), .ZN(n9342) );
  NAND2_X2 U13022 ( .A1(n9342), .A2(n6515), .ZN(n9740) );
  XNOR2_X2 U13023 ( .A(n12053), .B(n9342), .ZN(n9750) );
  MUX2_X2 U13024 ( .A(regBoiz_regfile_0__5_), .B(regBoiz_regfile_1__5_), .S(
        net369161), .Z(n9344) );
  MUX2_X2 U13025 ( .A(regBoiz_regfile_2__5_), .B(regBoiz_regfile_3__5_), .S(
        net369228), .Z(n9343) );
  MUX2_X2 U13026 ( .A(n9344), .B(n9343), .S(n6805), .Z(n9348) );
  MUX2_X2 U13027 ( .A(regBoiz_regfile_4__5_), .B(regBoiz_regfile_5__5_), .S(
        net369236), .Z(n9346) );
  MUX2_X2 U13028 ( .A(regBoiz_regfile_6__5_), .B(regBoiz_regfile_7__5_), .S(
        net369244), .Z(n9345) );
  MUX2_X2 U13029 ( .A(n9346), .B(n9345), .S(n6805), .Z(n9347) );
  MUX2_X2 U13030 ( .A(n9348), .B(n9347), .S(n6823), .Z(n9356) );
  MUX2_X2 U13031 ( .A(regBoiz_regfile_8__5_), .B(regBoiz_regfile_9__5_), .S(
        net377337), .Z(n9350) );
  MUX2_X2 U13032 ( .A(regBoiz_regfile_10__5_), .B(regBoiz_regfile_11__5_), .S(
        net369147), .Z(n9349) );
  MUX2_X2 U13033 ( .A(n9350), .B(n9349), .S(n6805), .Z(n9354) );
  MUX2_X2 U13034 ( .A(regBoiz_regfile_12__5_), .B(regBoiz_regfile_13__5_), .S(
        net378318), .Z(n9352) );
  MUX2_X2 U13035 ( .A(regBoiz_regfile_14__5_), .B(regBoiz_regfile_15__5_), .S(
        net369157), .Z(n9351) );
  MUX2_X2 U13036 ( .A(n9352), .B(n9351), .S(n6805), .Z(n9353) );
  MUX2_X2 U13037 ( .A(n9354), .B(n9353), .S(n6823), .Z(n9355) );
  MUX2_X2 U13038 ( .A(n9356), .B(n9355), .S(n6830), .Z(n9372) );
  MUX2_X2 U13039 ( .A(regBoiz_regfile_16__5_), .B(regBoiz_regfile_17__5_), .S(
        net369155), .Z(n9358) );
  MUX2_X2 U13040 ( .A(regBoiz_regfile_18__5_), .B(regBoiz_regfile_19__5_), .S(
        net369144), .Z(n9357) );
  MUX2_X2 U13041 ( .A(n9358), .B(n9357), .S(n6805), .Z(n9362) );
  MUX2_X2 U13042 ( .A(regBoiz_regfile_20__5_), .B(regBoiz_regfile_21__5_), .S(
        net369164), .Z(n9360) );
  MUX2_X2 U13043 ( .A(regBoiz_regfile_22__5_), .B(regBoiz_regfile_23__5_), .S(
        net369154), .Z(n9359) );
  MUX2_X2 U13044 ( .A(n9360), .B(n9359), .S(n6805), .Z(n9361) );
  MUX2_X2 U13045 ( .A(n9362), .B(n9361), .S(n6823), .Z(n9370) );
  MUX2_X2 U13046 ( .A(regBoiz_regfile_24__5_), .B(regBoiz_regfile_25__5_), .S(
        net369145), .Z(n9364) );
  MUX2_X2 U13047 ( .A(regBoiz_regfile_26__5_), .B(regBoiz_regfile_27__5_), .S(
        net369155), .Z(n9363) );
  MUX2_X2 U13048 ( .A(n9364), .B(n9363), .S(n6805), .Z(n9368) );
  MUX2_X2 U13049 ( .A(regBoiz_regfile_28__5_), .B(regBoiz_regfile_29__5_), .S(
        net369156), .Z(n9366) );
  MUX2_X2 U13050 ( .A(regBoiz_regfile_30__5_), .B(regBoiz_regfile_31__5_), .S(
        net369155), .Z(n9365) );
  MUX2_X2 U13051 ( .A(n9366), .B(n9365), .S(n6805), .Z(n9367) );
  MUX2_X2 U13052 ( .A(n9368), .B(n9367), .S(n6823), .Z(n9369) );
  MUX2_X2 U13053 ( .A(n9370), .B(n9369), .S(n6830), .Z(n9371) );
  MUX2_X2 U13054 ( .A(n9372), .B(n9371), .S(n6834), .Z(n13205) );
  NAND2_X2 U13055 ( .A1(n9718), .A2(n13205), .ZN(n9374) );
  NAND2_X2 U13056 ( .A1(daddr[26]), .A2(n6547), .ZN(n9373) );
  INV_X4 U13057 ( .A(n12309), .ZN(n9524) );
  XNOR2_X2 U13058 ( .A(n5762), .B(n9524), .ZN(n9375) );
  INV_X4 U13059 ( .A(n9375), .ZN(n9451) );
  INV_X4 U13060 ( .A(n9376), .ZN(n9379) );
  OAI21_X4 U13061 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(n9755) );
  MUX2_X2 U13062 ( .A(regBoiz_regfile_0__7_), .B(regBoiz_regfile_1__7_), .S(
        net369154), .Z(n9382) );
  MUX2_X2 U13063 ( .A(regBoiz_regfile_2__7_), .B(regBoiz_regfile_3__7_), .S(
        net369163), .Z(n9381) );
  MUX2_X2 U13064 ( .A(n9382), .B(n9381), .S(n6805), .Z(n9386) );
  MUX2_X2 U13065 ( .A(regBoiz_regfile_4__7_), .B(regBoiz_regfile_5__7_), .S(
        net369166), .Z(n9384) );
  MUX2_X2 U13066 ( .A(regBoiz_regfile_6__7_), .B(regBoiz_regfile_7__7_), .S(
        net369154), .Z(n9383) );
  MUX2_X2 U13067 ( .A(n9384), .B(n9383), .S(n6805), .Z(n9385) );
  MUX2_X2 U13068 ( .A(n9386), .B(n9385), .S(n6823), .Z(n9394) );
  MUX2_X2 U13069 ( .A(regBoiz_regfile_8__7_), .B(regBoiz_regfile_9__7_), .S(
        net369162), .Z(n9388) );
  MUX2_X2 U13070 ( .A(regBoiz_regfile_10__7_), .B(regBoiz_regfile_11__7_), .S(
        net369244), .Z(n9387) );
  MUX2_X2 U13071 ( .A(n9388), .B(n9387), .S(n6805), .Z(n9392) );
  MUX2_X2 U13072 ( .A(regBoiz_regfile_12__7_), .B(regBoiz_regfile_13__7_), .S(
        net369220), .Z(n9390) );
  MUX2_X2 U13073 ( .A(regBoiz_regfile_14__7_), .B(regBoiz_regfile_15__7_), .S(
        net378318), .Z(n9389) );
  MUX2_X2 U13074 ( .A(n9390), .B(n9389), .S(n6805), .Z(n9391) );
  MUX2_X2 U13075 ( .A(n9392), .B(n9391), .S(n6823), .Z(n9393) );
  MUX2_X2 U13076 ( .A(n9394), .B(n9393), .S(n6830), .Z(n9410) );
  MUX2_X2 U13077 ( .A(regBoiz_regfile_16__7_), .B(regBoiz_regfile_17__7_), .S(
        net369161), .Z(n9396) );
  MUX2_X2 U13078 ( .A(regBoiz_regfile_18__7_), .B(regBoiz_regfile_19__7_), .S(
        net377337), .Z(n9395) );
  MUX2_X2 U13079 ( .A(n9396), .B(n9395), .S(n6805), .Z(n9400) );
  MUX2_X2 U13080 ( .A(regBoiz_regfile_20__7_), .B(regBoiz_regfile_21__7_), .S(
        net369220), .Z(n9398) );
  MUX2_X2 U13081 ( .A(regBoiz_regfile_22__7_), .B(regBoiz_regfile_23__7_), .S(
        net369165), .Z(n9397) );
  MUX2_X2 U13082 ( .A(n9398), .B(n9397), .S(n6805), .Z(n9399) );
  MUX2_X2 U13083 ( .A(n9400), .B(n9399), .S(n6823), .Z(n9408) );
  MUX2_X2 U13084 ( .A(regBoiz_regfile_24__7_), .B(regBoiz_regfile_25__7_), .S(
        net369228), .Z(n9402) );
  MUX2_X2 U13085 ( .A(regBoiz_regfile_26__7_), .B(regBoiz_regfile_27__7_), .S(
        net369144), .Z(n9401) );
  MUX2_X2 U13086 ( .A(n9402), .B(n9401), .S(n6805), .Z(n9406) );
  MUX2_X2 U13087 ( .A(regBoiz_regfile_28__7_), .B(regBoiz_regfile_29__7_), .S(
        net369145), .Z(n9404) );
  MUX2_X2 U13088 ( .A(regBoiz_regfile_30__7_), .B(regBoiz_regfile_31__7_), .S(
        net369162), .Z(n9403) );
  MUX2_X2 U13089 ( .A(n9404), .B(n9403), .S(n6805), .Z(n9405) );
  MUX2_X2 U13090 ( .A(n9406), .B(n9405), .S(n6823), .Z(n9407) );
  MUX2_X2 U13091 ( .A(n9408), .B(n9407), .S(n6830), .Z(n9409) );
  MUX2_X2 U13092 ( .A(n9410), .B(n9409), .S(n6834), .Z(n13177) );
  NAND2_X2 U13093 ( .A1(n9718), .A2(n13177), .ZN(n9412) );
  NAND2_X2 U13094 ( .A1(daddr[24]), .A2(n6547), .ZN(n9411) );
  INV_X4 U13095 ( .A(n12208), .ZN(n9558) );
  XNOR2_X2 U13096 ( .A(n5762), .B(n9558), .ZN(n9413) );
  INV_X4 U13097 ( .A(n9413), .ZN(n9414) );
  XNOR2_X2 U13098 ( .A(n10101), .B(n9414), .ZN(n9756) );
  INV_X4 U13099 ( .A(n6517), .ZN(n10089) );
  MUX2_X2 U13100 ( .A(regBoiz_regfile_0__6_), .B(regBoiz_regfile_1__6_), .S(
        net369212), .Z(n9416) );
  MUX2_X2 U13101 ( .A(regBoiz_regfile_2__6_), .B(regBoiz_regfile_3__6_), .S(
        net369147), .Z(n9415) );
  MUX2_X2 U13102 ( .A(n9416), .B(n9415), .S(n6803), .Z(n9420) );
  MUX2_X2 U13103 ( .A(regBoiz_regfile_4__6_), .B(regBoiz_regfile_5__6_), .S(
        net369145), .Z(n9418) );
  MUX2_X2 U13104 ( .A(regBoiz_regfile_6__6_), .B(regBoiz_regfile_7__6_), .S(
        net369244), .Z(n9417) );
  MUX2_X2 U13105 ( .A(n9418), .B(n9417), .S(n6805), .Z(n9419) );
  MUX2_X2 U13106 ( .A(n9420), .B(n9419), .S(n6823), .Z(n9428) );
  MUX2_X2 U13107 ( .A(regBoiz_regfile_8__6_), .B(regBoiz_regfile_9__6_), .S(
        net378318), .Z(n9422) );
  MUX2_X2 U13108 ( .A(regBoiz_regfile_10__6_), .B(regBoiz_regfile_11__6_), .S(
        net377338), .Z(n9421) );
  MUX2_X2 U13109 ( .A(n9422), .B(n9421), .S(n6805), .Z(n9426) );
  MUX2_X2 U13110 ( .A(regBoiz_regfile_12__6_), .B(regBoiz_regfile_13__6_), .S(
        net369228), .Z(n9424) );
  MUX2_X2 U13111 ( .A(regBoiz_regfile_14__6_), .B(regBoiz_regfile_15__6_), .S(
        net369212), .Z(n9423) );
  MUX2_X2 U13112 ( .A(n9424), .B(n9423), .S(n6805), .Z(n9425) );
  MUX2_X2 U13113 ( .A(n9426), .B(n9425), .S(n6823), .Z(n9427) );
  MUX2_X2 U13114 ( .A(n9428), .B(n9427), .S(n6830), .Z(n9444) );
  MUX2_X2 U13115 ( .A(regBoiz_regfile_16__6_), .B(regBoiz_regfile_17__6_), .S(
        net369144), .Z(n9430) );
  MUX2_X2 U13116 ( .A(regBoiz_regfile_18__6_), .B(regBoiz_regfile_19__6_), .S(
        net369144), .Z(n9429) );
  MUX2_X2 U13117 ( .A(n9430), .B(n9429), .S(n6805), .Z(n9434) );
  MUX2_X2 U13118 ( .A(regBoiz_regfile_20__6_), .B(regBoiz_regfile_21__6_), .S(
        net369165), .Z(n9432) );
  MUX2_X2 U13119 ( .A(regBoiz_regfile_22__6_), .B(regBoiz_regfile_23__6_), .S(
        net369155), .Z(n9431) );
  MUX2_X2 U13120 ( .A(n9432), .B(n9431), .S(n6805), .Z(n9433) );
  MUX2_X2 U13121 ( .A(n9434), .B(n9433), .S(n6821), .Z(n9442) );
  MUX2_X2 U13122 ( .A(regBoiz_regfile_24__6_), .B(regBoiz_regfile_25__6_), .S(
        net369244), .Z(n9436) );
  MUX2_X2 U13123 ( .A(regBoiz_regfile_26__6_), .B(regBoiz_regfile_27__6_), .S(
        net369156), .Z(n9435) );
  MUX2_X2 U13124 ( .A(n9436), .B(n9435), .S(n6805), .Z(n9440) );
  MUX2_X2 U13125 ( .A(regBoiz_regfile_28__6_), .B(regBoiz_regfile_29__6_), .S(
        net369157), .Z(n9438) );
  MUX2_X2 U13126 ( .A(regBoiz_regfile_30__6_), .B(regBoiz_regfile_31__6_), .S(
        net369246), .Z(n9437) );
  MUX2_X2 U13127 ( .A(n9438), .B(n9437), .S(n6806), .Z(n9439) );
  MUX2_X2 U13128 ( .A(n9440), .B(n9439), .S(n6821), .Z(n9441) );
  MUX2_X2 U13129 ( .A(n9442), .B(n9441), .S(n6830), .Z(n9443) );
  MUX2_X2 U13130 ( .A(n9444), .B(n9443), .S(n6834), .Z(n13167) );
  NAND2_X2 U13131 ( .A1(n9718), .A2(n13167), .ZN(n9446) );
  NAND2_X2 U13132 ( .A1(daddr[25]), .A2(n6547), .ZN(n9445) );
  INV_X4 U13133 ( .A(n12207), .ZN(n9536) );
  XNOR2_X2 U13134 ( .A(n5762), .B(n9536), .ZN(n9447) );
  INV_X4 U13135 ( .A(n9447), .ZN(n9448) );
  XNOR2_X2 U13136 ( .A(n10089), .B(n9448), .ZN(n9767) );
  INV_X4 U13137 ( .A(n9767), .ZN(n9450) );
  NAND2_X2 U13138 ( .A1(n9448), .A2(n6517), .ZN(n9449) );
  OAI21_X4 U13139 ( .B1(n9768), .B2(n9450), .A(n9449), .ZN(n9735) );
  NAND3_X4 U13140 ( .A1(n9740), .A2(n9742), .A3(n9741), .ZN(n9454) );
  NAND3_X4 U13141 ( .A1(n9454), .A2(n9455), .A3(n9743), .ZN(n9745) );
  INV_X4 U13142 ( .A(n9460), .ZN(n9482) );
  XNOR2_X2 U13143 ( .A(n9462), .B(n9461), .ZN(n12941) );
  INV_X4 U13144 ( .A(n12941), .ZN(n9476) );
  XNOR2_X2 U13145 ( .A(n9468), .B(n9467), .ZN(n13071) );
  INV_X4 U13146 ( .A(n9470), .ZN(n9471) );
  XNOR2_X2 U13147 ( .A(n9472), .B(n9471), .ZN(n13059) );
  XNOR2_X2 U13148 ( .A(n9474), .B(n9473), .ZN(n13047) );
  INV_X4 U13149 ( .A(n9479), .ZN(n9480) );
  MUX2_X2 U13150 ( .A(n9722), .B(n5288), .S(n9486), .Z(n9487) );
  NAND2_X2 U13151 ( .A1(aluBoi_aluBoi_shft_srlout[21]), .A2(n5381), .ZN(n9490)
         );
  NAND2_X2 U13152 ( .A1(n9488), .A2(n10428), .ZN(n9489) );
  NAND3_X2 U13153 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(n13142) );
  MUX2_X2 U13154 ( .A(n9722), .B(n5288), .S(n9492), .Z(n9493) );
  MUX2_X2 U13155 ( .A(n9722), .B(n5288), .S(n9497), .Z(n9498) );
  NAND2_X2 U13156 ( .A1(aluBoi_aluBoi_shft_srlout[20]), .A2(n5381), .ZN(n9501)
         );
  NAND2_X2 U13157 ( .A1(n9499), .A2(n10427), .ZN(n9500) );
  NAND3_X2 U13158 ( .A1(n9502), .A2(n9501), .A3(n9500), .ZN(n13131) );
  MUX2_X2 U13159 ( .A(n9722), .B(n5288), .S(n9503), .Z(n9504) );
  NAND2_X2 U13160 ( .A1(aluBoi_aluBoi_shft_srlout[19]), .A2(n5381), .ZN(n9507)
         );
  NAND2_X2 U13161 ( .A1(n9505), .A2(n10423), .ZN(n9506) );
  NAND3_X2 U13162 ( .A1(n9508), .A2(n9507), .A3(n9506), .ZN(n13092) );
  INV_X4 U13163 ( .A(n13092), .ZN(n9522) );
  OAI21_X4 U13164 ( .B1(n6616), .B2(n6564), .A(n6561), .ZN(n9509) );
  NAND2_X2 U13165 ( .A1(n9509), .A2(n13525), .ZN(n9514) );
  NAND2_X2 U13166 ( .A1(aluBoi_aluBoi_shft_srlout[3]), .A2(n5381), .ZN(n9513)
         );
  INV_X4 U13167 ( .A(n13525), .ZN(n10372) );
  MUX2_X2 U13168 ( .A(n9680), .B(n6564), .S(n10372), .Z(n9510) );
  NAND2_X2 U13169 ( .A1(n9510), .A2(n6561), .ZN(n9511) );
  NAND2_X2 U13170 ( .A1(n9511), .A2(n6616), .ZN(n9512) );
  NAND3_X2 U13171 ( .A1(n9514), .A2(n9513), .A3(n9512), .ZN(n13250) );
  MUX2_X2 U13172 ( .A(n9722), .B(n5288), .S(n9515), .Z(n9516) );
  NAND2_X2 U13173 ( .A1(aluBoi_aluBoi_shft_srlout[18]), .A2(n6566), .ZN(n9519)
         );
  NAND2_X2 U13174 ( .A1(n9517), .A2(n10424), .ZN(n9518) );
  NAND3_X2 U13175 ( .A1(n9520), .A2(n9519), .A3(n9518), .ZN(n13102) );
  MUX2_X2 U13176 ( .A(n9722), .B(n5288), .S(n9524), .Z(n9525) );
  NAND2_X2 U13177 ( .A1(aluBoi_aluBoi_shft_srlout[26]), .A2(n6566), .ZN(n9528)
         );
  NAND2_X2 U13178 ( .A1(n9526), .A2(n12309), .ZN(n9527) );
  NAND3_X2 U13179 ( .A1(n9529), .A2(n9528), .A3(n9527), .ZN(n13209) );
  INV_X4 U13180 ( .A(n13209), .ZN(n9544) );
  MUX2_X2 U13181 ( .A(n9722), .B(n5288), .S(n9530), .Z(n9531) );
  OAI21_X4 U13182 ( .B1(n6562), .B2(n9531), .A(n6513), .ZN(n9535) );
  NAND2_X2 U13183 ( .A1(aluBoi_aluBoi_shft_srlout[28]), .A2(n6566), .ZN(n9534)
         );
  NAND2_X2 U13184 ( .A1(n9532), .A2(n12211), .ZN(n9533) );
  NAND3_X4 U13185 ( .A1(n9535), .A2(n9534), .A3(n9533), .ZN(n13191) );
  INV_X4 U13186 ( .A(n13191), .ZN(n9543) );
  MUX2_X2 U13187 ( .A(n9722), .B(n5288), .S(n9536), .Z(n9537) );
  NAND2_X2 U13188 ( .A1(aluBoi_aluBoi_shft_srlout[25]), .A2(n6566), .ZN(n9540)
         );
  OAI21_X4 U13189 ( .B1(n6517), .B2(n6564), .A(n6561), .ZN(n9538) );
  NAND2_X2 U13190 ( .A1(n9538), .A2(n12207), .ZN(n9539) );
  NAND3_X2 U13191 ( .A1(n9541), .A2(n9540), .A3(n9539), .ZN(n13171) );
  INV_X4 U13192 ( .A(n13171), .ZN(n9542) );
  MUX2_X2 U13193 ( .A(n9722), .B(n5288), .S(n9545), .Z(n9546) );
  NAND2_X2 U13194 ( .A1(aluBoi_aluBoi_shft_srlout[27]), .A2(n6566), .ZN(n9549)
         );
  OAI21_X4 U13195 ( .B1(n6515), .B2(n6564), .A(n6561), .ZN(n9547) );
  NAND2_X2 U13196 ( .A1(n9547), .A2(n10431), .ZN(n9548) );
  NAND3_X2 U13197 ( .A1(n9550), .A2(n9549), .A3(n9548), .ZN(n13199) );
  MUX2_X2 U13198 ( .A(n9722), .B(n5288), .S(n9551), .Z(n9552) );
  NAND2_X2 U13199 ( .A1(aluBoi_aluBoi_shft_srlout[22]), .A2(n6566), .ZN(n9555)
         );
  OAI21_X4 U13200 ( .B1(net368572), .B2(n6564), .A(n6561), .ZN(n9553) );
  NAND2_X2 U13201 ( .A1(n9553), .A2(n10429), .ZN(n9554) );
  NAND3_X2 U13202 ( .A1(n9556), .A2(n9555), .A3(n9554), .ZN(n13151) );
  MUX2_X2 U13203 ( .A(n9722), .B(n5288), .S(n9558), .Z(n9559) );
  NAND2_X2 U13204 ( .A1(aluBoi_aluBoi_shft_srlout[24]), .A2(n6566), .ZN(n9562)
         );
  NAND2_X2 U13205 ( .A1(n9560), .A2(n12208), .ZN(n9561) );
  NAND3_X2 U13206 ( .A1(n9563), .A2(n9562), .A3(n9561), .ZN(n13181) );
  NAND2_X2 U13207 ( .A1(n9564), .A2(n10430), .ZN(n9569) );
  NAND2_X2 U13208 ( .A1(aluBoi_aluBoi_shft_srlout[23]), .A2(n6566), .ZN(n9568)
         );
  MUX2_X2 U13209 ( .A(n9722), .B(n5288), .S(n9565), .Z(n9566) );
  NAND3_X2 U13210 ( .A1(n9569), .A2(n9568), .A3(n9567), .ZN(n13161) );
  OAI21_X4 U13211 ( .B1(n6614), .B2(n6564), .A(n6561), .ZN(n9570) );
  NAND2_X2 U13212 ( .A1(n9570), .A2(net376579), .ZN(n9575) );
  NAND2_X2 U13213 ( .A1(aluBoi_aluBoi_shft_srlout[2]), .A2(n6566), .ZN(n9574)
         );
  MUX2_X2 U13214 ( .A(n9680), .B(n6564), .S(net361801), .Z(n9571) );
  NAND2_X2 U13215 ( .A1(n9571), .A2(n6561), .ZN(n9572) );
  NAND2_X2 U13216 ( .A1(n9572), .A2(n6614), .ZN(n9573) );
  NAND3_X2 U13217 ( .A1(n9575), .A2(n9574), .A3(n9573), .ZN(n13259) );
  MUX2_X2 U13218 ( .A(n9722), .B(n5288), .S(n9576), .Z(n9577) );
  OAI21_X4 U13219 ( .B1(n6562), .B2(n9577), .A(n6509), .ZN(n9581) );
  NAND2_X2 U13220 ( .A1(aluBoi_aluBoi_shft_srlout[30]), .A2(n6566), .ZN(n9580)
         );
  NAND2_X2 U13221 ( .A1(n9578), .A2(n12312), .ZN(n9579) );
  NAND3_X4 U13222 ( .A1(n9581), .A2(n9580), .A3(n9579), .ZN(n13224) );
  OAI21_X4 U13223 ( .B1(n6606), .B2(n6563), .A(n6561), .ZN(n9582) );
  NAND2_X2 U13224 ( .A1(n9582), .A2(net368498), .ZN(n9587) );
  NAND2_X2 U13225 ( .A1(aluBoi_aluBoi_shft_srlout[1]), .A2(n6566), .ZN(n9586)
         );
  MUX2_X2 U13226 ( .A(n9680), .B(n6564), .S(net362224), .Z(n9583) );
  NAND2_X2 U13227 ( .A1(n9583), .A2(n6561), .ZN(n9584) );
  NAND2_X2 U13228 ( .A1(n9584), .A2(n6606), .ZN(n9585) );
  NAND3_X2 U13229 ( .A1(n9587), .A2(n9586), .A3(n9585), .ZN(n13270) );
  MUX2_X2 U13230 ( .A(n9722), .B(n5288), .S(n9588), .Z(n9589) );
  NAND2_X2 U13231 ( .A1(aluBoi_aluBoi_shft_srlout[16]), .A2(n6566), .ZN(n9592)
         );
  NAND2_X2 U13232 ( .A1(n9590), .A2(n10426), .ZN(n9591) );
  NAND3_X2 U13233 ( .A1(n9593), .A2(n9592), .A3(n9591), .ZN(n13124) );
  NAND2_X2 U13234 ( .A1(n9594), .A2(n12491), .ZN(n9599) );
  NAND2_X2 U13235 ( .A1(aluBoi_aluBoi_shft_srlout[29]), .A2(n6566), .ZN(n9598)
         );
  MUX2_X2 U13236 ( .A(n9722), .B(n5288), .S(n9595), .Z(n9596) );
  MUX2_X2 U13237 ( .A(n9722), .B(n5288), .S(n9600), .Z(n9601) );
  NAND2_X2 U13238 ( .A1(aluBoi_aluBoi_shft_srlout[17]), .A2(n6566), .ZN(n9604)
         );
  NAND2_X2 U13239 ( .A1(n9602), .A2(n10425), .ZN(n9603) );
  NAND3_X2 U13240 ( .A1(n9605), .A2(n9604), .A3(n9603), .ZN(n13113) );
  NAND4_X2 U13241 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n9645)
         );
  MUX2_X2 U13242 ( .A(n9722), .B(n5288), .S(n9610), .Z(n9611) );
  MUX2_X2 U13243 ( .A(n9722), .B(n5288), .S(n9615), .Z(n9616) );
  AOI22_X2 U13244 ( .A1(n9617), .A2(n10417), .B1(aluBoi_aluBoi_shft_srlout[10]), .B2(n5381), .ZN(n9618) );
  NAND2_X2 U13245 ( .A1(aluBoi_aluBoi_shft_srlout[4]), .A2(n5381), .ZN(n9623)
         );
  MUX2_X2 U13246 ( .A(n9722), .B(n5288), .S(net362485), .Z(n9621) );
  NAND3_X2 U13247 ( .A1(n9624), .A2(n9623), .A3(n9622), .ZN(n13012) );
  MUX2_X2 U13248 ( .A(n9722), .B(n5288), .S(n9625), .Z(n9626) );
  NAND2_X2 U13249 ( .A1(aluBoi_aluBoi_shft_srlout[8]), .A2(n6566), .ZN(n9629)
         );
  NAND2_X2 U13250 ( .A1(n9627), .A2(n10414), .ZN(n9628) );
  NAND3_X2 U13251 ( .A1(n9630), .A2(n9629), .A3(n9628), .ZN(n13020) );
  MUX2_X2 U13252 ( .A(n9722), .B(n5288), .S(n9631), .Z(n9632) );
  NOR2_X4 U13253 ( .A1(n6562), .A2(n9632), .ZN(n9636) );
  OAI21_X4 U13254 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n13031) );
  MUX2_X2 U13255 ( .A(n9722), .B(n5288), .S(n9637), .Z(n9638) );
  AOI22_X2 U13256 ( .A1(n9639), .A2(n10413), .B1(aluBoi_aluBoi_shft_srlout[9]), 
        .B2(n5381), .ZN(n9640) );
  NAND2_X2 U13257 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  NAND4_X2 U13258 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9777)
         );
  MUX2_X2 U13259 ( .A(n9722), .B(n5288), .S(n9651), .Z(n9652) );
  INV_X4 U13260 ( .A(n6539), .ZN(n9655) );
  AOI22_X2 U13261 ( .A1(n9653), .A2(n10421), .B1(aluBoi_aluBoi_shft_srlout[11]), .B2(n5381), .ZN(n9654) );
  MUX2_X2 U13262 ( .A(n9680), .B(n6564), .S(n9661), .Z(n9657) );
  AOI21_X2 U13263 ( .B1(aluBoi_aluBoi_shft_srlout[13]), .B2(n5381), .A(n9658), 
        .ZN(n9662) );
  INV_X4 U13264 ( .A(n9659), .ZN(n9660) );
  NAND2_X2 U13265 ( .A1(n9662), .A2(n5713), .ZN(n13061) );
  MUX2_X2 U13266 ( .A(n9680), .B(n6564), .S(n9664), .Z(n9663) );
  NAND2_X2 U13267 ( .A1(n9663), .A2(n6561), .ZN(n9669) );
  NAND2_X2 U13268 ( .A1(aluBoi_aluBoi_shft_srlout[12]), .A2(n6566), .ZN(n9666)
         );
  INV_X4 U13269 ( .A(n9666), .ZN(n9667) );
  AOI211_X4 U13270 ( .C1(n9669), .C2(n6384), .A(n9668), .B(n9667), .ZN(n13073)
         );
  MUX2_X2 U13271 ( .A(n9680), .B(n6564), .S(n9671), .Z(n9670) );
  NAND2_X2 U13272 ( .A1(n9670), .A2(n6561), .ZN(n9676) );
  NAND2_X2 U13273 ( .A1(n5288), .A2(n11067), .ZN(n9672) );
  NAND2_X2 U13274 ( .A1(aluBoi_aluBoi_shft_srlout[14]), .A2(n5381), .ZN(n9673)
         );
  INV_X4 U13275 ( .A(n9673), .ZN(n9674) );
  NAND2_X2 U13276 ( .A1(aluBoi_aluBoi_shft_srlout[0]), .A2(n6566), .ZN(n9687)
         );
  XNOR2_X2 U13277 ( .A(n9678), .B(n9677), .ZN(n9679) );
  NAND2_X2 U13278 ( .A1(n13220), .A2(n9679), .ZN(n9686) );
  MUX2_X2 U13279 ( .A(n9680), .B(n6563), .S(n6613), .Z(n9681) );
  NAND2_X2 U13280 ( .A1(n9681), .A2(n6561), .ZN(n9684) );
  NAND3_X2 U13281 ( .A1(n9687), .A2(n9686), .A3(n9685), .ZN(n13283) );
  MUX2_X2 U13282 ( .A(regBoiz_regfile_0__0_), .B(regBoiz_regfile_1__0_), .S(
        net369222), .Z(n9689) );
  MUX2_X2 U13283 ( .A(regBoiz_regfile_2__0_), .B(regBoiz_regfile_3__0_), .S(
        net369244), .Z(n9688) );
  MUX2_X2 U13284 ( .A(n9689), .B(n9688), .S(n6806), .Z(n9693) );
  MUX2_X2 U13285 ( .A(regBoiz_regfile_4__0_), .B(regBoiz_regfile_5__0_), .S(
        net377337), .Z(n9691) );
  MUX2_X2 U13286 ( .A(regBoiz_regfile_6__0_), .B(regBoiz_regfile_7__0_), .S(
        net369246), .Z(n9690) );
  MUX2_X2 U13287 ( .A(n9691), .B(n9690), .S(n6806), .Z(n9692) );
  MUX2_X2 U13288 ( .A(n9693), .B(n9692), .S(n6821), .Z(n9701) );
  MUX2_X2 U13289 ( .A(regBoiz_regfile_8__0_), .B(regBoiz_regfile_9__0_), .S(
        net369230), .Z(n9695) );
  MUX2_X2 U13290 ( .A(regBoiz_regfile_10__0_), .B(regBoiz_regfile_11__0_), .S(
        net378318), .Z(n9694) );
  MUX2_X2 U13291 ( .A(n9695), .B(n9694), .S(n6806), .Z(n9699) );
  MUX2_X2 U13292 ( .A(regBoiz_regfile_12__0_), .B(regBoiz_regfile_13__0_), .S(
        net369147), .Z(n9697) );
  MUX2_X2 U13293 ( .A(regBoiz_regfile_14__0_), .B(regBoiz_regfile_15__0_), .S(
        net369246), .Z(n9696) );
  MUX2_X2 U13294 ( .A(n9697), .B(n9696), .S(n6806), .Z(n9698) );
  MUX2_X2 U13295 ( .A(n9699), .B(n9698), .S(n6821), .Z(n9700) );
  MUX2_X2 U13296 ( .A(n9701), .B(n9700), .S(n6830), .Z(n9717) );
  MUX2_X2 U13297 ( .A(regBoiz_regfile_16__0_), .B(regBoiz_regfile_17__0_), .S(
        net378318), .Z(n9703) );
  MUX2_X2 U13298 ( .A(regBoiz_regfile_18__0_), .B(regBoiz_regfile_19__0_), .S(
        net369144), .Z(n9702) );
  MUX2_X2 U13299 ( .A(n9703), .B(n9702), .S(n6806), .Z(n9707) );
  MUX2_X2 U13300 ( .A(regBoiz_regfile_20__0_), .B(regBoiz_regfile_21__0_), .S(
        net378318), .Z(n9705) );
  MUX2_X2 U13301 ( .A(regBoiz_regfile_22__0_), .B(regBoiz_regfile_23__0_), .S(
        net369145), .Z(n9704) );
  MUX2_X2 U13302 ( .A(n9705), .B(n9704), .S(n6806), .Z(n9706) );
  MUX2_X2 U13303 ( .A(n9707), .B(n9706), .S(n6821), .Z(n9715) );
  MUX2_X2 U13304 ( .A(regBoiz_regfile_24__0_), .B(regBoiz_regfile_25__0_), .S(
        net369145), .Z(n9709) );
  MUX2_X2 U13305 ( .A(regBoiz_regfile_26__0_), .B(regBoiz_regfile_27__0_), .S(
        net378318), .Z(n9708) );
  MUX2_X2 U13306 ( .A(n9709), .B(n9708), .S(n6806), .Z(n9713) );
  MUX2_X2 U13307 ( .A(regBoiz_regfile_28__0_), .B(regBoiz_regfile_29__0_), .S(
        net369147), .Z(n9711) );
  MUX2_X2 U13308 ( .A(regBoiz_regfile_30__0_), .B(regBoiz_regfile_31__0_), .S(
        net369164), .Z(n9710) );
  MUX2_X2 U13309 ( .A(n9711), .B(n9710), .S(n6806), .Z(n9712) );
  MUX2_X2 U13310 ( .A(n9713), .B(n9712), .S(n6821), .Z(n9714) );
  MUX2_X2 U13311 ( .A(n9715), .B(n9714), .S(n6830), .Z(n9716) );
  MUX2_X2 U13312 ( .A(n9717), .B(n9716), .S(n6834), .Z(n13372) );
  NAND2_X2 U13313 ( .A1(n9718), .A2(n13372), .ZN(n9721) );
  NAND2_X2 U13314 ( .A1(n6547), .A2(daddr[31]), .ZN(n9720) );
  INV_X4 U13315 ( .A(n10497), .ZN(n9730) );
  MUX2_X2 U13316 ( .A(n9722), .B(n5288), .S(n9730), .Z(n9723) );
  NAND2_X2 U13317 ( .A1(n9724), .A2(n10497), .ZN(n9725) );
  NAND2_X2 U13318 ( .A1(n9726), .A2(n9725), .ZN(n13513) );
  INV_X4 U13319 ( .A(n6509), .ZN(n9729) );
  OAI21_X4 U13320 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9780) );
  XNOR2_X2 U13321 ( .A(n6565), .B(n9730), .ZN(n9778) );
  INV_X4 U13322 ( .A(n9778), .ZN(n9731) );
  XNOR2_X2 U13323 ( .A(n12183), .B(n9731), .ZN(n9779) );
  NAND2_X2 U13324 ( .A1(aluBoi_aluBoi_shft_sllout[31]), .A2(n12940), .ZN(
        n13509) );
  NAND2_X2 U13325 ( .A1(aluBoi_aluBoi_shft_srlout[31]), .A2(n5381), .ZN(n13511) );
  INV_X4 U13326 ( .A(n9781), .ZN(n9734) );
  NAND2_X2 U13327 ( .A1(aluBoi_aluBoi_shft_sraout[26]), .A2(n12944), .ZN(n9738) );
  NAND2_X2 U13328 ( .A1(aluBoi_aluBoi_shft_sllout[26]), .A2(n12940), .ZN(n9737) );
  INV_X4 U13329 ( .A(n9742), .ZN(n9744) );
  AND2_X2 U13330 ( .A1(aluBoi_aluBoi_shft_sraout[29]), .A2(n12944), .ZN(n9746)
         );
  AOI21_X2 U13331 ( .B1(aluBoi_aluBoi_shft_sllout[29]), .B2(n12940), .A(n9746), 
        .ZN(n9747) );
  INV_X4 U13332 ( .A(aluBoi_aluBoi_shft_sraout[27]), .ZN(n9754) );
  NAND2_X2 U13333 ( .A1(aluBoi_aluBoi_shft_sllout[27]), .A2(n12940), .ZN(n9752) );
  INV_X4 U13334 ( .A(aluBoi_aluBoi_shft_sllout[24]), .ZN(n9759) );
  NAND2_X2 U13335 ( .A1(aluBoi_aluBoi_shft_sraout[24]), .A2(n12944), .ZN(n9757) );
  INV_X4 U13336 ( .A(aluBoi_aluBoi_shft_sraout[28]), .ZN(n9765) );
  XNOR2_X2 U13337 ( .A(n9762), .B(n9761), .ZN(n9764) );
  NAND2_X2 U13338 ( .A1(aluBoi_aluBoi_shft_sllout[28]), .A2(n12940), .ZN(n9763) );
  NAND2_X2 U13339 ( .A1(aluBoi_aluBoi_shft_sraout[25]), .A2(n12944), .ZN(n9770) );
  NAND2_X2 U13340 ( .A1(aluBoi_aluBoi_shft_sllout[25]), .A2(n12940), .ZN(n9769) );
  OAI211_X2 U13341 ( .C1(n9771), .C2(n13222), .A(n9770), .B(n9769), .ZN(n13172) );
  NAND4_X2 U13342 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(n9776)
         );
  XNOR2_X2 U13343 ( .A(n9783), .B(n9782), .ZN(n2844) );
  INV_X4 U13344 ( .A(n2844), .ZN(n13575) );
  INV_X4 U13345 ( .A(ifInst[26]), .ZN(n13539) );
  NOR2_X4 U13346 ( .A1(n6511), .A2(n6509), .ZN(n9902) );
  NAND2_X2 U13347 ( .A1(n10562), .A2(net368548), .ZN(n10568) );
  OAI21_X4 U13348 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n10914) );
  NAND3_X2 U13349 ( .A1(n11726), .A2(n9804), .A3(n9803), .ZN(n9807) );
  NAND2_X2 U13350 ( .A1(n9805), .A2(n11769), .ZN(n9806) );
  NOR3_X4 U13351 ( .A1(n9809), .A2(n9810), .A3(n9811), .ZN(n9900) );
  INV_X4 U13352 ( .A(n9812), .ZN(n9817) );
  NOR2_X4 U13353 ( .A1(n9817), .A2(n9816), .ZN(n11477) );
  NAND2_X2 U13354 ( .A1(n9818), .A2(net367045), .ZN(n9821) );
  NAND3_X2 U13355 ( .A1(n9821), .A2(n9820), .A3(n6787), .ZN(n9827) );
  NOR2_X4 U13356 ( .A1(n11054), .A2(n9823), .ZN(n9824) );
  NAND3_X4 U13357 ( .A1(n9827), .A2(n9826), .A3(net362297), .ZN(n9828) );
  INV_X4 U13358 ( .A(n11180), .ZN(n9837) );
  INV_X4 U13359 ( .A(n9833), .ZN(n9836) );
  INV_X4 U13360 ( .A(n9834), .ZN(n9835) );
  INV_X4 U13361 ( .A(n9846), .ZN(n9852) );
  INV_X4 U13362 ( .A(n9854), .ZN(n9860) );
  NAND3_X2 U13363 ( .A1(n9857), .A2(n9856), .A3(n9855), .ZN(n9858) );
  INV_X4 U13364 ( .A(n9858), .ZN(n9859) );
  AOI21_X4 U13365 ( .B1(n7750), .B2(n9860), .A(n9859), .ZN(n9865) );
  INV_X4 U13366 ( .A(n9862), .ZN(n9863) );
  NAND2_X2 U13367 ( .A1(n9865), .A2(n9864), .ZN(n9873) );
  NAND3_X2 U13368 ( .A1(n9867), .A2(n9866), .A3(net375506), .ZN(n9868) );
  INV_X4 U13369 ( .A(n9868), .ZN(n9871) );
  OAI21_X4 U13370 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(n10779) );
  NAND2_X2 U13371 ( .A1(n9875), .A2(net368548), .ZN(n10778) );
  INV_X4 U13372 ( .A(net363049), .ZN(net363046) );
  OAI21_X4 U13373 ( .B1(net363046), .B2(net363047), .A(n9876), .ZN(n11181) );
  INV_X4 U13374 ( .A(n9885), .ZN(n9886) );
  NAND3_X4 U13375 ( .A1(n6066), .A2(n9887), .A3(n9886), .ZN(n10697) );
  INV_X4 U13376 ( .A(n9888), .ZN(n9891) );
  NAND2_X2 U13377 ( .A1(n9888), .A2(net368548), .ZN(n9889) );
  OAI21_X4 U13378 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n11192) );
  INV_X4 U13379 ( .A(n11183), .ZN(n9896) );
  NAND3_X4 U13380 ( .A1(n11244), .A2(n11243), .A3(n11245), .ZN(n11722) );
  NOR2_X4 U13381 ( .A1(n9903), .A2(n5556), .ZN(n9904) );
  NAND2_X2 U13382 ( .A1(ifInst[27]), .A2(ifInst[26]), .ZN(n13426) );
  INV_X4 U13383 ( .A(ifInst[28]), .ZN(n13493) );
  INV_X4 U13384 ( .A(ifInst[27]), .ZN(n13491) );
  OAI21_X4 U13385 ( .B1(n13426), .B2(n13324), .A(n12917), .ZN(n9905) );
  INV_X4 U13386 ( .A(ifInst[29]), .ZN(n13495) );
  NAND2_X2 U13387 ( .A1(n9905), .A2(n13495), .ZN(n12916) );
  NOR2_X4 U13388 ( .A1(aluifJRflag), .A2(n12916), .ZN(n9906) );
  NAND3_X4 U13389 ( .A1(n9940), .A2(n6239), .A3(n9906), .ZN(n9988) );
  NAND2_X2 U13390 ( .A1(ifOut_94_), .A2(ifInst[25]), .ZN(n9938) );
  XNOR2_X2 U13391 ( .A(ifOut_90_), .B(n5313), .ZN(n10073) );
  XNOR2_X2 U13392 ( .A(ifOut_89_), .B(ifInst[25]), .ZN(n10084) );
  XNOR2_X2 U13393 ( .A(ifOut_87_), .B(ifInst[23]), .ZN(n10112) );
  XNOR2_X2 U13394 ( .A(ifOut_85_), .B(ifInst[21]), .ZN(n10137) );
  XNOR2_X2 U13395 ( .A(ifOut_83_), .B(ifInst[19]), .ZN(n10166) );
  XNOR2_X2 U13396 ( .A(ifOut_81_), .B(ifInst[17]), .ZN(n10192) );
  XNOR2_X2 U13397 ( .A(ifOut_79_), .B(ifInst[15]), .ZN(n10220) );
  XNOR2_X2 U13398 ( .A(ifOut_77_), .B(ifInst[13]), .ZN(n10245) );
  XNOR2_X2 U13399 ( .A(ifOut_75_), .B(ifInst[11]), .ZN(n10270) );
  XNOR2_X2 U13400 ( .A(ifOut_73_), .B(ifInst[9]), .ZN(n10292) );
  XNOR2_X2 U13401 ( .A(ifOut_71_), .B(ifInst[7]), .ZN(n10324) );
  XNOR2_X2 U13402 ( .A(ifOut_69_), .B(ifInst[5]), .ZN(n10347) );
  XNOR2_X2 U13403 ( .A(ifOut_67_), .B(ifInst[3]), .ZN(n10376) );
  XNOR2_X2 U13404 ( .A(ifOut_65_), .B(idBoi_temPC_1_), .ZN(n10396) );
  INV_X4 U13405 ( .A(n10384), .ZN(n9908) );
  NAND2_X2 U13406 ( .A1(ifOut_67_), .A2(ifInst[3]), .ZN(n9909) );
  OAI21_X4 U13407 ( .B1(n10376), .B2(n10377), .A(n9909), .ZN(n10358) );
  XNOR2_X2 U13408 ( .A(ifOut_68_), .B(ifInst[4]), .ZN(n10357) );
  INV_X4 U13409 ( .A(n10357), .ZN(n9910) );
  NAND2_X2 U13410 ( .A1(ifOut_69_), .A2(ifInst[5]), .ZN(n9911) );
  XNOR2_X2 U13411 ( .A(ifOut_70_), .B(ifInst[6]), .ZN(n10338) );
  INV_X4 U13412 ( .A(n10338), .ZN(n9912) );
  NAND2_X2 U13413 ( .A1(ifOut_71_), .A2(ifInst[7]), .ZN(n9913) );
  OAI21_X4 U13414 ( .B1(n10324), .B2(n10325), .A(n9913), .ZN(n10306) );
  XNOR2_X2 U13415 ( .A(ifOut_72_), .B(ifInst[8]), .ZN(n10305) );
  INV_X4 U13416 ( .A(n10305), .ZN(n9914) );
  NAND2_X2 U13417 ( .A1(ifOut_73_), .A2(ifInst[9]), .ZN(n9915) );
  XNOR2_X2 U13418 ( .A(ifOut_74_), .B(ifInst[10]), .ZN(n10277) );
  INV_X4 U13419 ( .A(n10277), .ZN(n9916) );
  NAND2_X2 U13420 ( .A1(ifOut_75_), .A2(ifInst[11]), .ZN(n9917) );
  OAI21_X4 U13421 ( .B1(n10270), .B2(n10271), .A(n9917), .ZN(n10253) );
  XNOR2_X2 U13422 ( .A(ifOut_76_), .B(ifInst[12]), .ZN(n10252) );
  INV_X4 U13423 ( .A(n10252), .ZN(n9918) );
  NAND2_X2 U13424 ( .A1(ifOut_77_), .A2(ifInst[13]), .ZN(n9919) );
  OAI21_X4 U13425 ( .B1(n10245), .B2(n10246), .A(n9919), .ZN(n10228) );
  XNOR2_X2 U13426 ( .A(ifOut_78_), .B(ifInst[14]), .ZN(n10227) );
  INV_X4 U13427 ( .A(n10227), .ZN(n9920) );
  NAND2_X2 U13428 ( .A1(ifOut_79_), .A2(ifInst[15]), .ZN(n9921) );
  OAI21_X4 U13429 ( .B1(n10220), .B2(n10221), .A(n9921), .ZN(n10210) );
  XNOR2_X2 U13430 ( .A(ifOut_80_), .B(ifInst[16]), .ZN(n10209) );
  INV_X4 U13431 ( .A(n10209), .ZN(n9922) );
  NAND2_X2 U13432 ( .A1(ifOut_81_), .A2(ifInst[17]), .ZN(n9923) );
  XNOR2_X2 U13433 ( .A(ifOut_82_), .B(ifInst[18]), .ZN(n10173) );
  INV_X4 U13434 ( .A(n10173), .ZN(n9924) );
  NAND2_X2 U13435 ( .A1(ifOut_83_), .A2(ifInst[19]), .ZN(n9925) );
  XNOR2_X2 U13436 ( .A(ifOut_84_), .B(ifInst[20]), .ZN(n10149) );
  INV_X4 U13437 ( .A(n10149), .ZN(n9926) );
  NAND2_X2 U13438 ( .A1(ifOut_85_), .A2(ifInst[21]), .ZN(n9927) );
  OAI21_X4 U13439 ( .B1(n10138), .B2(n10137), .A(n9927), .ZN(n10126) );
  XNOR2_X2 U13440 ( .A(ifOut_86_), .B(ifInst[22]), .ZN(n10125) );
  INV_X4 U13441 ( .A(n10125), .ZN(n9928) );
  NAND2_X2 U13442 ( .A1(ifOut_87_), .A2(ifInst[23]), .ZN(n9929) );
  OAI21_X4 U13443 ( .B1(n10113), .B2(n10112), .A(n9929), .ZN(n10100) );
  NAND2_X2 U13444 ( .A1(ifOut_89_), .A2(n5313), .ZN(n9930) );
  OAI21_X4 U13445 ( .B1(n10085), .B2(n10084), .A(n9930), .ZN(n10074) );
  INV_X4 U13446 ( .A(n10074), .ZN(n9932) );
  NAND2_X2 U13447 ( .A1(ifOut_90_), .A2(n5313), .ZN(n9931) );
  OAI21_X4 U13448 ( .B1(n10073), .B2(n9932), .A(n9931), .ZN(n10057) );
  XNOR2_X2 U13449 ( .A(ifOut_91_), .B(ifInst[25]), .ZN(n10058) );
  INV_X4 U13450 ( .A(n10058), .ZN(n9933) );
  NAND2_X2 U13451 ( .A1(n10057), .A2(n9933), .ZN(n9934) );
  INV_X4 U13452 ( .A(n9934), .ZN(n10047) );
  AOI211_X4 U13453 ( .C1(ifOut_92_), .C2(ifInst[25]), .A(n10047), .B(n5351), 
        .ZN(n9937) );
  OAI22_X2 U13454 ( .A1(ifOut_93_), .A2(ifInst[25]), .B1(ifOut_92_), .B2(
        ifInst[25]), .ZN(n9936) );
  NAND2_X2 U13455 ( .A1(ifOut_93_), .A2(ifInst[25]), .ZN(n9935) );
  OAI21_X4 U13456 ( .B1(n9937), .B2(n9936), .A(n9935), .ZN(n9939) );
  NAND4_X2 U13457 ( .A1(ifOut_95_), .A2(ifInst[25]), .A3(n9938), .A4(n10001), 
        .ZN(n9946) );
  INV_X4 U13458 ( .A(ifInst[25]), .ZN(n13488) );
  NAND3_X4 U13459 ( .A1(n10001), .A2(ifInst[25]), .A3(n5461), .ZN(n10000) );
  NAND2_X2 U13460 ( .A1(n13301), .A2(ifInst[27]), .ZN(n13427) );
  INV_X4 U13461 ( .A(n13427), .ZN(n13321) );
  INV_X4 U13462 ( .A(n9994), .ZN(n9943) );
  INV_X4 U13463 ( .A(n9942), .ZN(n9995) );
  NAND3_X4 U13464 ( .A1(n9943), .A2(n6548), .A3(n9995), .ZN(n10139) );
  AOI21_X4 U13465 ( .B1(n9944), .B2(n10000), .A(n10139), .ZN(n9945) );
  XNOR2_X2 U13466 ( .A(n6569), .B(n5517), .ZN(n10060) );
  XNOR2_X2 U13467 ( .A(n6568), .B(n5516), .ZN(n10086) );
  XNOR2_X2 U13468 ( .A(n6568), .B(n5514), .ZN(n10127) );
  XNOR2_X2 U13469 ( .A(n6568), .B(n5513), .ZN(n10151) );
  XNOR2_X2 U13470 ( .A(n6568), .B(n5518), .ZN(n10164) );
  XNOR2_X2 U13471 ( .A(n6568), .B(n5486), .ZN(n10175) );
  XNOR2_X2 U13472 ( .A(n6568), .B(n5523), .ZN(n10190) );
  NAND2_X2 U13473 ( .A1(idOut_100_), .A2(aluBoi_imm32w_14_), .ZN(n10203) );
  XNOR2_X2 U13474 ( .A(idOut_99_), .B(aluBoi_imm32w_13_), .ZN(n10242) );
  XNOR2_X2 U13475 ( .A(idOut_97_), .B(aluBoi_imm32w_11_), .ZN(n10267) );
  XNOR2_X2 U13476 ( .A(idOut_95_), .B(aluBoi_imm32w_9_), .ZN(n10296) );
  XNOR2_X2 U13477 ( .A(idOut_93_), .B(aluBoi_imm32w_7_), .ZN(n10321) );
  XNOR2_X2 U13478 ( .A(idOut_91_), .B(aluBoi_imm32w_5_), .ZN(n10350) );
  XNOR2_X2 U13479 ( .A(idOut_89_), .B(aluBoi_imm32w_3_), .ZN(n10373) );
  NOR2_X4 U13480 ( .A1(idOut_87_), .A2(aluBoi_imm32w_1_), .ZN(n9949) );
  NAND2_X2 U13481 ( .A1(idOut_87_), .A2(aluBoi_imm32w_1_), .ZN(n9948) );
  OAI21_X4 U13482 ( .B1(n9949), .B2(n10392), .A(n9948), .ZN(n10387) );
  NAND2_X2 U13483 ( .A1(idOut_89_), .A2(aluBoi_imm32w_3_), .ZN(n9950) );
  OAI21_X4 U13484 ( .B1(n10374), .B2(n10373), .A(n9950), .ZN(n10360) );
  XNOR2_X2 U13485 ( .A(idOut_90_), .B(aluBoi_imm32w_4_), .ZN(n10359) );
  INV_X4 U13486 ( .A(n10359), .ZN(n9951) );
  NAND2_X2 U13487 ( .A1(idOut_91_), .A2(aluBoi_imm32w_5_), .ZN(n9952) );
  OAI21_X4 U13488 ( .B1(n10351), .B2(n10350), .A(n9952), .ZN(n10337) );
  XNOR2_X2 U13489 ( .A(idOut_92_), .B(aluBoi_imm32w_6_), .ZN(n10336) );
  INV_X4 U13490 ( .A(n10336), .ZN(n9953) );
  NAND2_X2 U13491 ( .A1(idOut_93_), .A2(aluBoi_imm32w_7_), .ZN(n9954) );
  OAI21_X4 U13492 ( .B1(n10322), .B2(n10321), .A(n9954), .ZN(n10308) );
  XNOR2_X2 U13493 ( .A(idOut_94_), .B(aluBoi_imm32w_8_), .ZN(n10307) );
  INV_X4 U13494 ( .A(n10307), .ZN(n9955) );
  NAND2_X2 U13495 ( .A1(idOut_95_), .A2(aluBoi_imm32w_9_), .ZN(n9956) );
  OAI21_X4 U13496 ( .B1(n10295), .B2(n10296), .A(n9956), .ZN(n10280) );
  XNOR2_X2 U13497 ( .A(idOut_96_), .B(aluBoi_imm32w_10_), .ZN(n10279) );
  INV_X4 U13498 ( .A(n10279), .ZN(n9957) );
  NAND2_X2 U13499 ( .A1(idOut_97_), .A2(aluBoi_imm32w_11_), .ZN(n9958) );
  OAI21_X4 U13500 ( .B1(n10268), .B2(n10267), .A(n9958), .ZN(n10255) );
  XNOR2_X2 U13501 ( .A(idOut_98_), .B(aluBoi_imm32w_12_), .ZN(n10254) );
  INV_X4 U13502 ( .A(n10254), .ZN(n9959) );
  NAND2_X2 U13503 ( .A1(idOut_99_), .A2(aluBoi_imm32w_13_), .ZN(n9960) );
  OAI21_X4 U13504 ( .B1(n10243), .B2(n10242), .A(n9960), .ZN(n10230) );
  XNOR2_X2 U13505 ( .A(idOut_100_), .B(aluBoi_imm32w_14_), .ZN(n10229) );
  INV_X4 U13506 ( .A(n10229), .ZN(n9961) );
  NAND2_X2 U13507 ( .A1(n10230), .A2(n9961), .ZN(n10202) );
  NAND2_X2 U13508 ( .A1(idOut_101_), .A2(aluBoi_imm32w_15_), .ZN(n10204) );
  NAND3_X2 U13509 ( .A1(n10203), .A2(n10202), .A3(n10204), .ZN(n9964) );
  XNOR2_X2 U13510 ( .A(idOut_101_), .B(aluBoi_imm32w_15_), .ZN(n10218) );
  NAND2_X2 U13511 ( .A1(n10218), .A2(n10204), .ZN(n9963) );
  XNOR2_X2 U13512 ( .A(n6568), .B(n5512), .ZN(n9962) );
  INV_X4 U13513 ( .A(n9962), .ZN(n10208) );
  NAND3_X2 U13514 ( .A1(n9964), .A2(n9963), .A3(n10208), .ZN(n9965) );
  NOR2_X4 U13515 ( .A1(n5750), .A2(n10151), .ZN(n9967) );
  NOR2_X4 U13516 ( .A1(n9967), .A2(n9966), .ZN(n10135) );
  XNOR2_X2 U13517 ( .A(n6568), .B(n5504), .ZN(n10134) );
  NOR2_X4 U13518 ( .A1(n10127), .A2(n9968), .ZN(n9970) );
  NOR2_X4 U13519 ( .A1(n9970), .A2(n9969), .ZN(n10111) );
  XNOR2_X2 U13520 ( .A(n6568), .B(n5515), .ZN(n10110) );
  NOR2_X4 U13521 ( .A1(n10111), .A2(n10110), .ZN(n9972) );
  NOR2_X4 U13522 ( .A1(n9972), .A2(n9971), .ZN(n10099) );
  XNOR2_X2 U13523 ( .A(n6568), .B(n5524), .ZN(n10098) );
  NOR2_X4 U13524 ( .A1(n5915), .A2(n10086), .ZN(n9974) );
  NOR2_X4 U13525 ( .A1(n9974), .A2(n9973), .ZN(n10072) );
  XNOR2_X2 U13526 ( .A(n6569), .B(n5505), .ZN(n10071) );
  NOR2_X4 U13527 ( .A1(n10060), .A2(n9975), .ZN(n9977) );
  NAND2_X2 U13528 ( .A1(idOut_115_), .A2(idOut_114_), .ZN(n9978) );
  INV_X4 U13529 ( .A(n9982), .ZN(n10005) );
  MUX2_X2 U13530 ( .A(n6569), .B(n5349), .S(n10005), .Z(n9985) );
  NAND2_X2 U13531 ( .A1(idOut_116_), .A2(n6569), .ZN(n9981) );
  OAI211_X2 U13532 ( .C1(n9982), .C2(n9981), .A(n10008), .B(n5554), .ZN(n9983)
         );
  INV_X4 U13533 ( .A(n12830), .ZN(n10299) );
  NAND2_X2 U13534 ( .A1(n10299), .A2(iaddr[9]), .ZN(n10285) );
  INV_X4 U13535 ( .A(n10285), .ZN(n12599) );
  INV_X4 U13536 ( .A(n12876), .ZN(n12840) );
  NAND2_X2 U13537 ( .A1(n12599), .A2(n5347), .ZN(n12826) );
  INV_X4 U13538 ( .A(n12826), .ZN(n10284) );
  NAND2_X2 U13539 ( .A1(n10284), .A2(iaddr[10]), .ZN(n12810) );
  INV_X4 U13540 ( .A(n12810), .ZN(n10264) );
  NAND2_X2 U13541 ( .A1(n10264), .A2(iaddr[11]), .ZN(n12811) );
  INV_X4 U13542 ( .A(n12811), .ZN(n10259) );
  INV_X4 U13543 ( .A(n12786), .ZN(n10215) );
  NAND2_X2 U13544 ( .A1(iaddr[15]), .A2(n10215), .ZN(n12770) );
  INV_X4 U13545 ( .A(n12770), .ZN(n10199) );
  NAND2_X2 U13546 ( .A1(iaddr[16]), .A2(n10199), .ZN(n12765) );
  INV_X4 U13547 ( .A(n12765), .ZN(n10186) );
  NAND2_X2 U13548 ( .A1(iaddr[17]), .A2(n10186), .ZN(n12750) );
  INV_X4 U13549 ( .A(n12750), .ZN(n10181) );
  NAND2_X2 U13550 ( .A1(iaddr[18]), .A2(n10181), .ZN(n12745) );
  INV_X4 U13551 ( .A(n12745), .ZN(n10161) );
  INV_X4 U13552 ( .A(n12730), .ZN(n10156) );
  NAND2_X2 U13553 ( .A1(iaddr[20]), .A2(n10156), .ZN(n12725) );
  INV_X4 U13554 ( .A(n12725), .ZN(n10144) );
  INV_X4 U13555 ( .A(n12710), .ZN(n10122) );
  NAND2_X2 U13556 ( .A1(iaddr[22]), .A2(n10122), .ZN(n12705) );
  INV_X4 U13557 ( .A(n12705), .ZN(n9986) );
  NOR2_X4 U13558 ( .A1(n12687), .A2(n5559), .ZN(n12667) );
  NAND2_X2 U13559 ( .A1(iaddr[27]), .A2(n5886), .ZN(n12645) );
  INV_X4 U13560 ( .A(n12645), .ZN(n9987) );
  INV_X4 U13561 ( .A(n12613), .ZN(n9989) );
  NAND2_X2 U13562 ( .A1(n9989), .A2(n10369), .ZN(n9991) );
  MUX2_X2 U13563 ( .A(n9991), .B(n9990), .S(iaddr[31]), .Z(n9997) );
  INV_X4 U13564 ( .A(n9992), .ZN(difHold) );
  NAND3_X4 U13565 ( .A1(n9995), .A2(n9994), .A3(n9993), .ZN(n10403) );
  NAND4_X2 U13566 ( .A1(n9999), .A2(n9998), .A3(n9997), .A4(n9996), .ZN(n4558)
         );
  INV_X4 U13567 ( .A(n10000), .ZN(n10004) );
  XNOR2_X2 U13568 ( .A(ifOut_94_), .B(ifInst[25]), .ZN(n10002) );
  MUX2_X2 U13569 ( .A(n10002), .B(n5557), .S(n10001), .Z(n10003) );
  NAND2_X2 U13570 ( .A1(idOut_116_), .A2(n6569), .ZN(n10007) );
  XNOR2_X2 U13571 ( .A(idOut_116_), .B(n6569), .ZN(n10006) );
  MUX2_X2 U13572 ( .A(n10007), .B(n10006), .S(n10005), .Z(n10009) );
  AOI21_X4 U13573 ( .B1(n10009), .B2(n10008), .A(n6577), .ZN(n10015) );
  NAND2_X2 U13574 ( .A1(n10369), .A2(n10010), .ZN(n10012) );
  MUX2_X2 U13575 ( .A(n10012), .B(n10011), .S(iaddr[30]), .Z(n10013) );
  NAND2_X2 U13576 ( .A1(n10013), .A2(n5712), .ZN(n10014) );
  NOR2_X4 U13577 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  NAND2_X2 U13578 ( .A1(n10017), .A2(n10016), .ZN(n4563) );
  NOR2_X4 U13579 ( .A1(n10047), .A2(n5351), .ZN(n10021) );
  INV_X4 U13580 ( .A(n10021), .ZN(n10018) );
  NAND2_X2 U13581 ( .A1(n10018), .A2(n13488), .ZN(n10020) );
  INV_X4 U13582 ( .A(n10020), .ZN(n10019) );
  NAND2_X2 U13583 ( .A1(n10021), .A2(ifInst[25]), .ZN(n10023) );
  INV_X4 U13584 ( .A(n10023), .ZN(n10024) );
  NAND4_X2 U13585 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10042) );
  MUX2_X2 U13586 ( .A(idOut_114_), .B(n5916), .S(n5017), .Z(n10029) );
  AOI21_X4 U13587 ( .B1(n5686), .B2(n10029), .A(n5350), .ZN(n10034) );
  INV_X4 U13588 ( .A(n10030), .ZN(n10031) );
  MUX2_X2 U13589 ( .A(n10032), .B(n10031), .S(n5916), .Z(n10033) );
  OAI21_X4 U13590 ( .B1(n10034), .B2(n10033), .A(n6576), .ZN(n10041) );
  MUX2_X2 U13591 ( .A(n10037), .B(n10036), .S(iaddr[29]), .Z(n10038) );
  NOR2_X4 U13592 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  NAND3_X4 U13593 ( .A1(n10041), .A2(n10042), .A3(n10040), .ZN(n4568) );
  XNOR2_X2 U13594 ( .A(n6568), .B(n5462), .ZN(n10044) );
  NOR2_X4 U13595 ( .A1(ifOut_91_), .A2(n10047), .ZN(n10046) );
  MUX2_X2 U13596 ( .A(n10047), .B(n10046), .S(ifInst[25]), .Z(n10048) );
  XNOR2_X2 U13597 ( .A(ifOut_92_), .B(n10048), .ZN(n10055) );
  INV_X4 U13598 ( .A(n6513), .ZN(n12054) );
  NAND2_X2 U13599 ( .A1(n10049), .A2(n6548), .ZN(n10050) );
  MUX2_X2 U13600 ( .A(n10051), .B(n10050), .S(iaddr[28]), .Z(n10052) );
  OAI221_X2 U13601 ( .B1(n10056), .B2(n6577), .C1(n10055), .C2(n10139), .A(
        n10054), .ZN(n4573) );
  INV_X4 U13602 ( .A(n10057), .ZN(n10059) );
  XNOR2_X2 U13603 ( .A(n10059), .B(n10058), .ZN(n10070) );
  NAND2_X2 U13604 ( .A1(n6576), .A2(n10062), .ZN(n10069) );
  NOR2_X4 U13605 ( .A1(n12660), .A2(n6551), .ZN(n10065) );
  NAND2_X2 U13606 ( .A1(n6571), .A2(n12660), .ZN(n10063) );
  NAND2_X2 U13607 ( .A1(n10063), .A2(n6548), .ZN(n10064) );
  MUX2_X2 U13608 ( .A(n10065), .B(n10064), .S(iaddr[27]), .Z(n10066) );
  OAI211_X2 U13609 ( .C1(n10070), .C2(n10139), .A(n10069), .B(n10068), .ZN(
        n4578) );
  XNOR2_X2 U13610 ( .A(n10072), .B(n10071), .ZN(n10083) );
  INV_X4 U13611 ( .A(n10073), .ZN(n10075) );
  XNOR2_X2 U13612 ( .A(n10075), .B(n10074), .ZN(n10082) );
  NAND2_X2 U13613 ( .A1(n6571), .A2(n12666), .ZN(n10076) );
  NAND2_X2 U13614 ( .A1(n10076), .A2(n6548), .ZN(n10077) );
  MUX2_X2 U13615 ( .A(n10078), .B(n10077), .S(iaddr[26]), .Z(n10079) );
  OAI221_X2 U13616 ( .B1(n10083), .B2(n6577), .C1(n10082), .C2(n10139), .A(
        n10081), .ZN(n4583) );
  XNOR2_X2 U13617 ( .A(n10087), .B(n10086), .ZN(n10088) );
  NAND2_X2 U13618 ( .A1(n6576), .A2(n10088), .ZN(n10096) );
  INV_X4 U13619 ( .A(n12667), .ZN(n12681) );
  NAND2_X2 U13620 ( .A1(n6571), .A2(n12681), .ZN(n10090) );
  NAND2_X2 U13621 ( .A1(n10090), .A2(n6548), .ZN(n10091) );
  MUX2_X2 U13622 ( .A(n10092), .B(n10091), .S(iaddr[25]), .Z(n10093) );
  OAI211_X2 U13623 ( .C1(n10097), .C2(n10139), .A(n10096), .B(n10095), .ZN(
        n4588) );
  XNOR2_X2 U13624 ( .A(n10099), .B(n10098), .ZN(n10109) );
  XNOR2_X2 U13625 ( .A(n5352), .B(n10100), .ZN(n10108) );
  NAND2_X2 U13626 ( .A1(n10102), .A2(n6548), .ZN(n10103) );
  MUX2_X2 U13627 ( .A(n10104), .B(n10103), .S(iaddr[24]), .Z(n10105) );
  NOR2_X4 U13628 ( .A1(n10106), .A2(n10105), .ZN(n10107) );
  OAI221_X2 U13629 ( .B1(n10109), .B2(n6577), .C1(n10108), .C2(n10139), .A(
        n10107), .ZN(n4593) );
  XNOR2_X2 U13630 ( .A(n10111), .B(n10110), .ZN(n10121) );
  NOR2_X4 U13631 ( .A1(net360550), .A2(n6573), .ZN(n10118) );
  NAND2_X2 U13632 ( .A1(n10114), .A2(n6548), .ZN(n10115) );
  MUX2_X2 U13633 ( .A(n10116), .B(n10115), .S(iaddr[23]), .Z(n10117) );
  NOR2_X4 U13634 ( .A1(n10118), .A2(n10117), .ZN(n10119) );
  OAI221_X2 U13635 ( .B1(n10121), .B2(n6577), .C1(n10120), .C2(n10139), .A(
        n10119), .ZN(n4598) );
  NAND2_X2 U13636 ( .A1(n6575), .A2(net368572), .ZN(n10133) );
  NAND2_X2 U13637 ( .A1(n10369), .A2(n10122), .ZN(n10124) );
  MUX2_X2 U13638 ( .A(n10124), .B(n10123), .S(iaddr[22]), .Z(n10132) );
  XNOR2_X2 U13639 ( .A(n10126), .B(n10125), .ZN(n10130) );
  AOI22_X2 U13640 ( .A1(n10408), .A2(n10130), .B1(n6576), .B2(n10129), .ZN(
        n10131) );
  NOR2_X4 U13641 ( .A1(n11524), .A2(n6573), .ZN(n10143) );
  XNOR2_X2 U13642 ( .A(n10135), .B(n10134), .ZN(n10136) );
  NOR3_X4 U13643 ( .A1(n10143), .A2(n10142), .A3(n10141), .ZN(n10148) );
  NAND2_X2 U13644 ( .A1(n10369), .A2(n10144), .ZN(n10146) );
  MUX2_X2 U13645 ( .A(n10146), .B(n10145), .S(iaddr[21]), .Z(n10147) );
  NAND2_X2 U13646 ( .A1(n10148), .A2(n10147), .ZN(n4608) );
  XNOR2_X2 U13647 ( .A(n10150), .B(n10149), .ZN(n10155) );
  AOI221_X2 U13648 ( .B1(n10408), .B2(n10155), .C1(n6576), .C2(n10154), .A(
        n10153), .ZN(n10160) );
  NAND2_X2 U13649 ( .A1(n10369), .A2(n10156), .ZN(n10158) );
  MUX2_X2 U13650 ( .A(n10158), .B(n10157), .S(iaddr[20]), .Z(n10159) );
  NAND2_X2 U13651 ( .A1(n10160), .A2(n10159), .ZN(n4613) );
  NAND2_X2 U13652 ( .A1(n10369), .A2(n10161), .ZN(n10163) );
  MUX2_X2 U13653 ( .A(n10163), .B(n10162), .S(iaddr[19]), .Z(n10172) );
  INV_X4 U13654 ( .A(n10166), .ZN(n10168) );
  AOI22_X2 U13655 ( .A1(n6576), .A2(n10170), .B1(n10408), .B2(n10169), .ZN(
        n10171) );
  NAND3_X2 U13656 ( .A1(n10172), .A2(n5710), .A3(n10171), .ZN(n4618) );
  XNOR2_X2 U13657 ( .A(n10174), .B(n10173), .ZN(n10180) );
  AOI221_X2 U13658 ( .B1(n10408), .B2(n10180), .C1(n6576), .C2(n10179), .A(
        n10178), .ZN(n10185) );
  NAND2_X2 U13659 ( .A1(n10369), .A2(n10181), .ZN(n10183) );
  MUX2_X2 U13660 ( .A(n10183), .B(n10182), .S(iaddr[18]), .Z(n10184) );
  NAND2_X2 U13661 ( .A1(n10185), .A2(n10184), .ZN(n4623) );
  NAND2_X2 U13662 ( .A1(n10369), .A2(n10186), .ZN(n10188) );
  MUX2_X2 U13663 ( .A(n10188), .B(n10187), .S(iaddr[17]), .Z(n10198) );
  XNOR2_X2 U13664 ( .A(n10191), .B(n10190), .ZN(n10196) );
  INV_X4 U13665 ( .A(n10192), .ZN(n10194) );
  AOI22_X2 U13666 ( .A1(n6576), .A2(n10196), .B1(n10408), .B2(n10195), .ZN(
        n10197) );
  NAND3_X2 U13667 ( .A1(n10198), .A2(n5704), .A3(n10197), .ZN(n4628) );
  NAND2_X2 U13668 ( .A1(n10369), .A2(n10199), .ZN(n10201) );
  MUX2_X2 U13669 ( .A(n10201), .B(n10200), .S(iaddr[16]), .Z(n10214) );
  NAND2_X2 U13670 ( .A1(n10203), .A2(n10202), .ZN(n10219) );
  INV_X4 U13671 ( .A(n10218), .ZN(n10206) );
  INV_X4 U13672 ( .A(n10204), .ZN(n10205) );
  AOI21_X4 U13673 ( .B1(n10219), .B2(n10206), .A(n10205), .ZN(n10207) );
  XNOR2_X2 U13674 ( .A(n10208), .B(n10207), .ZN(n10212) );
  XNOR2_X2 U13675 ( .A(n10210), .B(n10209), .ZN(n10211) );
  AOI22_X2 U13676 ( .A1(n6576), .A2(n10212), .B1(n10408), .B2(n10211), .ZN(
        n10213) );
  NAND3_X2 U13677 ( .A1(n10214), .A2(n5705), .A3(n10213), .ZN(n4633) );
  NAND2_X2 U13678 ( .A1(n10369), .A2(n10215), .ZN(n10217) );
  MUX2_X2 U13679 ( .A(n10217), .B(n10216), .S(iaddr[15]), .Z(n10226) );
  XNOR2_X2 U13680 ( .A(n10219), .B(n10218), .ZN(n10224) );
  INV_X4 U13681 ( .A(n10220), .ZN(n10222) );
  AOI22_X2 U13682 ( .A1(n6576), .A2(n10224), .B1(n10408), .B2(n10223), .ZN(
        n10225) );
  NAND3_X2 U13683 ( .A1(n10226), .A2(n5701), .A3(n10225), .ZN(n4638) );
  XNOR2_X2 U13684 ( .A(n10228), .B(n10227), .ZN(n10233) );
  XNOR2_X2 U13685 ( .A(n10230), .B(n10229), .ZN(n10232) );
  AOI221_X2 U13686 ( .B1(n10408), .B2(n10233), .C1(n6576), .C2(n10232), .A(
        n10231), .ZN(n10238) );
  NAND2_X2 U13687 ( .A1(n10369), .A2(n10234), .ZN(n10236) );
  MUX2_X2 U13688 ( .A(n10236), .B(n10235), .S(iaddr[14]), .Z(n10237) );
  NAND2_X2 U13689 ( .A1(n10238), .A2(n10237), .ZN(n4643) );
  NAND2_X2 U13690 ( .A1(n10369), .A2(n10239), .ZN(n10241) );
  MUX2_X2 U13691 ( .A(n10241), .B(n10240), .S(iaddr[13]), .Z(n10251) );
  INV_X4 U13692 ( .A(n10242), .ZN(n10244) );
  INV_X4 U13693 ( .A(n10245), .ZN(n10247) );
  AOI22_X2 U13694 ( .A1(n6576), .A2(n10249), .B1(n10408), .B2(n10248), .ZN(
        n10250) );
  NAND3_X2 U13695 ( .A1(n10251), .A2(n5706), .A3(n10250), .ZN(n4648) );
  XNOR2_X2 U13696 ( .A(n10253), .B(n10252), .ZN(n10258) );
  AOI221_X2 U13697 ( .B1(n10408), .B2(n10258), .C1(n6576), .C2(n10257), .A(
        n10256), .ZN(n10263) );
  NAND2_X2 U13698 ( .A1(n10369), .A2(n10259), .ZN(n10261) );
  MUX2_X2 U13699 ( .A(n10261), .B(n10260), .S(iaddr[12]), .Z(n10262) );
  NAND2_X2 U13700 ( .A1(n10263), .A2(n10262), .ZN(n4653) );
  NAND2_X2 U13701 ( .A1(n10369), .A2(n10264), .ZN(n10266) );
  MUX2_X2 U13702 ( .A(n10266), .B(n10265), .S(iaddr[11]), .Z(n10276) );
  INV_X4 U13703 ( .A(n10267), .ZN(n10269) );
  INV_X4 U13704 ( .A(n10270), .ZN(n10272) );
  AOI22_X2 U13705 ( .A1(n6576), .A2(n10274), .B1(n10408), .B2(n10273), .ZN(
        n10275) );
  NAND3_X2 U13706 ( .A1(n10276), .A2(n5707), .A3(n10275), .ZN(n4658) );
  XNOR2_X2 U13707 ( .A(n10278), .B(n10277), .ZN(n10283) );
  AOI221_X2 U13708 ( .B1(n10408), .B2(n10283), .C1(n6576), .C2(n10282), .A(
        n10281), .ZN(n10290) );
  NAND2_X2 U13709 ( .A1(n10369), .A2(n10284), .ZN(n10288) );
  MUX2_X2 U13710 ( .A(n10288), .B(n10287), .S(iaddr[10]), .Z(n10289) );
  NAND2_X2 U13711 ( .A1(n10290), .A2(n10289), .ZN(n4663) );
  AOI21_X4 U13712 ( .B1(n10408), .B2(n10294), .A(n10293), .ZN(n10304) );
  NAND2_X2 U13713 ( .A1(n6576), .A2(n10297), .ZN(n10303) );
  INV_X4 U13714 ( .A(n10344), .ZN(n10298) );
  NAND2_X2 U13715 ( .A1(n10299), .A2(n5647), .ZN(n12833) );
  NAND2_X2 U13716 ( .A1(n10369), .A2(n5347), .ZN(n10345) );
  NAND3_X4 U13717 ( .A1(n10304), .A2(n10303), .A3(n10302), .ZN(n4668) );
  XNOR2_X2 U13718 ( .A(n10306), .B(n10305), .ZN(n10312) );
  AOI221_X2 U13719 ( .B1(n10408), .B2(n10312), .C1(n6576), .C2(n10311), .A(
        n10310), .ZN(n10317) );
  NAND2_X2 U13720 ( .A1(n5347), .A2(iaddr[5]), .ZN(n12870) );
  INV_X4 U13721 ( .A(n12870), .ZN(n10331) );
  INV_X4 U13722 ( .A(n12853), .ZN(n10318) );
  INV_X4 U13723 ( .A(n12854), .ZN(n10313) );
  NAND2_X2 U13724 ( .A1(n10313), .A2(n10369), .ZN(n10315) );
  MUX2_X2 U13725 ( .A(n10315), .B(n10314), .S(iaddr[8]), .Z(n10316) );
  NAND2_X2 U13726 ( .A1(n10317), .A2(n10316), .ZN(n4673) );
  NAND2_X2 U13727 ( .A1(n10369), .A2(n10318), .ZN(n10320) );
  MUX2_X2 U13728 ( .A(n10320), .B(n10319), .S(iaddr[7]), .Z(n10330) );
  INV_X4 U13729 ( .A(n6541), .ZN(n10708) );
  INV_X4 U13730 ( .A(n10321), .ZN(n10323) );
  INV_X4 U13731 ( .A(n10324), .ZN(n10326) );
  AOI22_X2 U13732 ( .A1(n6576), .A2(n10328), .B1(n10408), .B2(n10327), .ZN(
        n10329) );
  NAND3_X2 U13733 ( .A1(n10330), .A2(n5708), .A3(n10329), .ZN(n4678) );
  NAND2_X2 U13734 ( .A1(n10369), .A2(n10331), .ZN(n10335) );
  MUX2_X2 U13735 ( .A(n10335), .B(n10334), .S(iaddr[6]), .Z(n10343) );
  INV_X4 U13736 ( .A(n6543), .ZN(n10575) );
  XNOR2_X2 U13737 ( .A(n10339), .B(n10338), .ZN(n10340) );
  AOI22_X2 U13738 ( .A1(n6576), .A2(n10341), .B1(n10408), .B2(n10340), .ZN(
        n10342) );
  NAND3_X2 U13739 ( .A1(n10343), .A2(n5709), .A3(n10342), .ZN(n4683) );
  MUX2_X2 U13740 ( .A(n10345), .B(n10298), .S(iaddr[5]), .Z(n10356) );
  INV_X4 U13741 ( .A(n10347), .ZN(n10349) );
  INV_X4 U13742 ( .A(n10350), .ZN(n10352) );
  AOI22_X2 U13743 ( .A1(n10408), .A2(n10354), .B1(n6576), .B2(n10353), .ZN(
        n10355) );
  NAND3_X2 U13744 ( .A1(n10356), .A2(n5703), .A3(n10355), .ZN(n4688) );
  XNOR2_X2 U13745 ( .A(n10358), .B(n10357), .ZN(n10363) );
  AOI221_X2 U13746 ( .B1(n10408), .B2(n10363), .C1(n6576), .C2(n10362), .A(
        n10361), .ZN(n10368) );
  INV_X4 U13747 ( .A(n12883), .ZN(n10364) );
  NAND2_X2 U13748 ( .A1(n10364), .A2(n10369), .ZN(n10366) );
  MUX2_X2 U13749 ( .A(n10366), .B(n10365), .S(iaddr[4]), .Z(n10367) );
  NAND2_X2 U13750 ( .A1(n10368), .A2(n10367), .ZN(n4693) );
  NAND2_X2 U13751 ( .A1(n10369), .A2(iaddr[2]), .ZN(n10371) );
  MUX2_X2 U13752 ( .A(n10371), .B(n10370), .S(iaddr[3]), .Z(n10382) );
  INV_X4 U13753 ( .A(n10376), .ZN(n10378) );
  AOI22_X2 U13754 ( .A1(n6576), .A2(n10380), .B1(n10408), .B2(n10379), .ZN(
        n10381) );
  NAND3_X2 U13755 ( .A1(n10382), .A2(n5702), .A3(n10381), .ZN(n4698) );
  MUX2_X2 U13756 ( .A(n6551), .B(n6548), .S(iaddr[2]), .Z(n10391) );
  AOI22_X2 U13757 ( .A1(n10408), .A2(n10389), .B1(n6576), .B2(n10388), .ZN(
        n10390) );
  NAND3_X2 U13758 ( .A1(n10391), .A2(n5711), .A3(n10390), .ZN(n4703) );
  INV_X4 U13759 ( .A(n10392), .ZN(n10393) );
  XNOR2_X2 U13760 ( .A(n10394), .B(n10393), .ZN(n10395) );
  NAND2_X2 U13761 ( .A1(n6576), .A2(n10395), .ZN(n10402) );
  NAND2_X2 U13762 ( .A1(n6575), .A2(net368498), .ZN(n10401) );
  NAND2_X2 U13763 ( .A1(iaddr[1]), .A2(n5390), .ZN(n10400) );
  NAND2_X2 U13764 ( .A1(n10408), .A2(n10398), .ZN(n10399) );
  NAND4_X2 U13765 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n4708) );
  NAND2_X2 U13766 ( .A1(iaddr[0]), .A2(n5390), .ZN(n10410) );
  NAND2_X2 U13767 ( .A1(n10408), .A2(n10407), .ZN(n10409) );
  MUX2_X2 U13768 ( .A(aluBoi_multBoi_temppp[2]), .B(n6606), .S(net367631), .Z(
        n13704) );
  MUX2_X2 U13769 ( .A(aluBoi_multBoi_temppp[6]), .B(n5020), .S(net368481), .Z(
        n13703) );
  MUX2_X2 U13770 ( .A(aluBoi_multBoi_temppp[10]), .B(n10413), .S(net368481), 
        .Z(n13696) );
  MUX2_X2 U13771 ( .A(aluBoi_multBoi_temppp[1]), .B(n6612), .S(net368481), .Z(
        n13702) );
  MUX2_X2 U13772 ( .A(aluBoi_multBoi_temppp[5]), .B(n6618), .S(net368481), .Z(
        n13701) );
  MUX2_X2 U13773 ( .A(aluBoi_multBoi_temppp[9]), .B(n10414), .S(net368481), 
        .Z(n13695) );
  MUX2_X2 U13774 ( .A(aluBoi_multBoi_temppp[4]), .B(n6616), .S(net368481), .Z(
        n13700) );
  MUX2_X2 U13775 ( .A(aluBoi_multBoi_temppp[8]), .B(n10415), .S(net367631), 
        .Z(n13694) );
  MUX2_X2 U13776 ( .A(aluBoi_multBoi_temppp[3]), .B(n6614), .S(net367631), .Z(
        n13699) );
  MUX2_X2 U13777 ( .A(aluBoi_multBoi_temppp[7]), .B(n10416), .S(net367631), 
        .Z(n13698) );
  MUX2_X2 U13778 ( .A(aluBoi_multBoi_temppp[11]), .B(n10417), .S(net367631), 
        .Z(n13697) );
  MUX2_X2 U13779 ( .A(aluBoi_multBoi_temppp[15]), .B(n10418), .S(net367631), 
        .Z(n13691) );
  MUX2_X2 U13780 ( .A(aluBoi_multBoi_temppp[14]), .B(n10419), .S(net367631), 
        .Z(n13690) );
  MUX2_X2 U13781 ( .A(aluBoi_multBoi_temppp[13]), .B(n10420), .S(net367631), 
        .Z(n13689) );
  MUX2_X2 U13782 ( .A(aluBoi_multBoi_temppp[12]), .B(n10421), .S(net367631), 
        .Z(n13693) );
  MUX2_X2 U13783 ( .A(aluBoi_multBoi_temppp[16]), .B(n10422), .S(net367631), 
        .Z(n13692) );
  MUX2_X2 U13784 ( .A(aluBoi_multBoi_temppp[20]), .B(n10423), .S(net367631), 
        .Z(n13685) );
  MUX2_X2 U13785 ( .A(aluBoi_multBoi_temppp[19]), .B(n10424), .S(net367631), 
        .Z(n13686) );
  MUX2_X2 U13786 ( .A(aluBoi_multBoi_temppp[18]), .B(n10425), .S(net367631), 
        .Z(n13687) );
  MUX2_X2 U13787 ( .A(aluBoi_multBoi_temppp[17]), .B(n10426), .S(net367631), 
        .Z(n13688) );
  MUX2_X2 U13788 ( .A(aluBoi_multBoi_temppp[21]), .B(n10427), .S(net367631), 
        .Z(n13682) );
  MUX2_X2 U13789 ( .A(aluBoi_multBoi_temppp[22]), .B(n10428), .S(net367631), 
        .Z(n13683) );
  MUX2_X2 U13790 ( .A(aluBoi_multBoi_temppp[23]), .B(n10429), .S(net367631), 
        .Z(n13680) );
  MUX2_X2 U13791 ( .A(aluBoi_multBoi_temppp[24]), .B(n10430), .S(net367631), 
        .Z(n13684) );
  MUX2_X2 U13792 ( .A(aluBoi_multBoi_temppp[28]), .B(n10431), .S(net367631), 
        .Z(aluBoi_multBoi_N34) );
  MUX2_X2 U13793 ( .A(n10446), .B(net362387), .S(net366927), .Z(n10447) );
  NAND2_X2 U13794 ( .A1(n6531), .A2(n10447), .ZN(n10448) );
  NOR2_X4 U13795 ( .A1(n10452), .A2(net368209), .ZN(n10456) );
  AOI21_X4 U13796 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(n10460) );
  AOI21_X4 U13797 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(n10465) );
  INV_X4 U13798 ( .A(n10466), .ZN(n10461) );
  NOR2_X4 U13799 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  XNOR2_X2 U13800 ( .A(n10465), .B(n10464), .ZN(net362317) );
  XNOR2_X2 U13801 ( .A(net362224), .B(net362256), .ZN(net362105) );
  INV_X4 U13802 ( .A(net362362), .ZN(net362361) );
  NAND2_X2 U13803 ( .A1(n10467), .A2(net362224), .ZN(n10473) );
  NAND2_X2 U13804 ( .A1(n10489), .A2(n10488), .ZN(net362218) );
  NAND2_X2 U13805 ( .A1(net368462), .A2(net375435), .ZN(n10470) );
  NAND2_X2 U13806 ( .A1(n10470), .A2(net345751), .ZN(n10491) );
  INV_X4 U13807 ( .A(n10491), .ZN(n10471) );
  OAI22_X2 U13808 ( .A1(net364246), .A2(net368467), .B1(net362105), .B2(
        net368211), .ZN(n10492) );
  NAND2_X2 U13809 ( .A1(net360904), .A2(n6251), .ZN(n10472) );
  NAND2_X2 U13810 ( .A1(n10474), .A2(net361801), .ZN(net362330) );
  OAI21_X4 U13811 ( .B1(n10481), .B2(n10480), .A(net362341), .ZN(n10482) );
  INV_X4 U13812 ( .A(n10483), .ZN(n10485) );
  XNOR2_X2 U13813 ( .A(n10486), .B(net362327), .ZN(net362134) );
  INV_X4 U13814 ( .A(net362318), .ZN(net362229) );
  NAND2_X2 U13815 ( .A1(net362229), .A2(net362230), .ZN(net362052) );
  NAND2_X2 U13816 ( .A1(n10489), .A2(n10488), .ZN(net362049) );
  AOI21_X4 U13817 ( .B1(net368444), .B2(net368185), .A(net362287), .ZN(
        net362311) );
  INV_X4 U13818 ( .A(net362016), .ZN(net362314) );
  AOI21_X4 U13819 ( .B1(net368436), .B2(net368179), .A(net362287), .ZN(n10654)
         );
  XNOR2_X2 U13820 ( .A(net362314), .B(n10654), .ZN(n10661) );
  XNOR2_X2 U13821 ( .A(n10661), .B(n5679), .ZN(n10662) );
  INV_X4 U13822 ( .A(n10490), .ZN(n10495) );
  XNOR2_X2 U13823 ( .A(aluBoi_multBoi_temppp[31]), .B(n10495), .ZN(n12311) );
  XNOR2_X2 U13824 ( .A(n10493), .B(n5678), .ZN(n12490) );
  NAND2_X2 U13825 ( .A1(net368467), .A2(net368211), .ZN(n12209) );
  NAND3_X4 U13826 ( .A1(aluBoi_multBoi_temppp[29]), .A2(net345751), .A3(n12209), .ZN(n12489) );
  INV_X4 U13827 ( .A(n12489), .ZN(n10494) );
  AOI22_X2 U13828 ( .A1(n12490), .A2(n10494), .B1(aluBoi_multBoi_temppp[30]), 
        .B2(n10493), .ZN(n12310) );
  NAND2_X2 U13829 ( .A1(aluBoi_multBoi_temppp[31]), .A2(n10495), .ZN(n10496)
         );
  OAI21_X4 U13830 ( .B1(n12311), .B2(n12310), .A(n10496), .ZN(n10663) );
  XOR2_X2 U13831 ( .A(n10662), .B(n10663), .Z(n10498) );
  MUX2_X2 U13832 ( .A(n10498), .B(n10497), .S(net367631), .Z(
        aluBoi_multBoi_N38) );
  INV_X4 U13833 ( .A(n10573), .ZN(n10607) );
  XNOR2_X2 U13834 ( .A(n10499), .B(n11230), .ZN(n10580) );
  OAI22_X2 U13835 ( .A1(n10500), .A2(net368436), .B1(n10580), .B2(net368179), 
        .ZN(n10599) );
  INV_X4 U13836 ( .A(n10599), .ZN(n10648) );
  NAND2_X2 U13837 ( .A1(net360821), .A2(n6545), .ZN(n10556) );
  INV_X4 U13838 ( .A(n10556), .ZN(n10517) );
  INV_X4 U13839 ( .A(n10502), .ZN(n10608) );
  INV_X4 U13840 ( .A(n10562), .ZN(n10504) );
  XNOR2_X2 U13841 ( .A(n10507), .B(n10506), .ZN(n10557) );
  NAND2_X2 U13842 ( .A1(net361984), .A2(n5310), .ZN(n10548) );
  NAND3_X4 U13843 ( .A1(n10518), .A2(net361801), .A3(net361802), .ZN(n10644)
         );
  NAND2_X2 U13844 ( .A1(net368201), .A2(n10644), .ZN(n10514) );
  INV_X4 U13845 ( .A(n10526), .ZN(n10530) );
  XNOR2_X2 U13846 ( .A(net362246), .B(n10531), .ZN(n10532) );
  INV_X4 U13847 ( .A(net362211), .ZN(net362223) );
  NAND2_X2 U13848 ( .A1(net362158), .A2(net362159), .ZN(n10541) );
  NAND3_X2 U13849 ( .A1(net362050), .A2(net362218), .A3(n10541), .ZN(n10542)
         );
  NAND2_X2 U13850 ( .A1(net360904), .A2(n6545), .ZN(n10637) );
  XNOR2_X2 U13851 ( .A(n10565), .B(n10564), .ZN(n10636) );
  NAND2_X2 U13852 ( .A1(net361802), .A2(net361801), .ZN(n10566) );
  INV_X4 U13853 ( .A(n10566), .ZN(n10721) );
  NAND3_X4 U13854 ( .A1(n10682), .A2(net361984), .A3(n5952), .ZN(n10725) );
  INV_X4 U13855 ( .A(n13523), .ZN(n10571) );
  INV_X4 U13856 ( .A(n10614), .ZN(n10572) );
  XNOR2_X2 U13857 ( .A(n10627), .B(n10577), .ZN(net361949) );
  INV_X4 U13858 ( .A(net361891), .ZN(net362125) );
  OAI22_X2 U13859 ( .A1(n10581), .A2(net368447), .B1(n10580), .B2(net368185), 
        .ZN(n10587) );
  OAI21_X4 U13860 ( .B1(net362156), .B2(net362157), .A(net362049), .ZN(n10583)
         );
  OAI211_X2 U13861 ( .C1(n10584), .C2(net377576), .A(net362053), .B(net362050), 
        .ZN(n10588) );
  INV_X4 U13862 ( .A(net362142), .ZN(net362127) );
  INV_X4 U13863 ( .A(net362092), .ZN(net362126) );
  NAND2_X2 U13864 ( .A1(net362096), .A2(net362097), .ZN(n10650) );
  OAI22_X2 U13865 ( .A1(net364246), .A2(net368436), .B1(n6441), .B2(net368179), 
        .ZN(n10594) );
  INV_X4 U13866 ( .A(n10594), .ZN(n10593) );
  XNOR2_X2 U13867 ( .A(n5743), .B(n10593), .ZN(n10655) );
  NAND3_X4 U13868 ( .A1(n10655), .A2(net362016), .A3(n10654), .ZN(n10657) );
  NAND3_X4 U13869 ( .A1(n10650), .A2(n10657), .A3(n10649), .ZN(n10596) );
  AOI21_X4 U13870 ( .B1(n10648), .B2(n10598), .A(n10597), .ZN(n10602) );
  INV_X4 U13871 ( .A(net362096), .ZN(net362095) );
  XNOR2_X2 U13872 ( .A(net362094), .B(net362095), .ZN(n10670) );
  NAND2_X2 U13873 ( .A1(net361891), .A2(net362092), .ZN(n10603) );
  NAND2_X2 U13874 ( .A1(net362091), .A2(n10603), .ZN(n10646) );
  XNOR2_X2 U13875 ( .A(net362194), .B(n5951), .ZN(net361889) );
  NAND2_X2 U13876 ( .A1(n10603), .A2(net378422), .ZN(n10604) );
  INV_X4 U13877 ( .A(n10604), .ZN(n10754) );
  NAND2_X2 U13878 ( .A1(n6541), .A2(n10684), .ZN(n10611) );
  NAND2_X2 U13879 ( .A1(n10616), .A2(n10615), .ZN(n10624) );
  NAND2_X2 U13880 ( .A1(n10714), .A2(n10625), .ZN(n10618) );
  NAND2_X2 U13881 ( .A1(n10620), .A2(n10619), .ZN(n10749) );
  INV_X4 U13882 ( .A(n10624), .ZN(n10626) );
  OAI21_X4 U13883 ( .B1(n10627), .B2(n10626), .A(n10625), .ZN(n10629) );
  OAI21_X4 U13884 ( .B1(n10628), .B2(net362053), .A(n10838), .ZN(n10643) );
  INV_X4 U13885 ( .A(n10630), .ZN(n10642) );
  XNOR2_X2 U13886 ( .A(n10633), .B(n10632), .ZN(n10842) );
  XNOR2_X2 U13887 ( .A(n10638), .B(n10639), .ZN(n10840) );
  NAND3_X4 U13888 ( .A1(n10643), .A2(n10642), .A3(n10641), .ZN(net361903) );
  NAND3_X4 U13889 ( .A1(n10749), .A2(net361903), .A3(n10750), .ZN(net361906)
         );
  XNOR2_X2 U13890 ( .A(n10644), .B(n6545), .ZN(n10759) );
  NAND2_X2 U13891 ( .A1(net359752), .A2(n6545), .ZN(n10645) );
  OAI21_X4 U13892 ( .B1(n10759), .B2(net368185), .A(n10645), .ZN(net361907) );
  XNOR2_X2 U13893 ( .A(net361906), .B(net361907), .ZN(net361827) );
  OAI22_X2 U13894 ( .A1(net362485), .A2(net368436), .B1(net368181), .B2(
        net362028), .ZN(net361893) );
  XNOR2_X2 U13895 ( .A(n10754), .B(net362026), .ZN(n10862) );
  XNOR2_X2 U13896 ( .A(n10871), .B(n5687), .ZN(n10868) );
  INV_X4 U13897 ( .A(n10646), .ZN(n10647) );
  XNOR2_X2 U13898 ( .A(n10648), .B(n10647), .ZN(n10672) );
  INV_X4 U13899 ( .A(n10672), .ZN(n10652) );
  XNOR2_X2 U13900 ( .A(n10652), .B(n10673), .ZN(n12314) );
  INV_X4 U13901 ( .A(n12314), .ZN(n10653) );
  NAND2_X2 U13902 ( .A1(aluBoi_multBoi_temppp[35]), .A2(n10653), .ZN(n10869)
         );
  NAND2_X2 U13903 ( .A1(n10654), .A2(net362016), .ZN(n10656) );
  NAND2_X2 U13904 ( .A1(n10656), .A2(n5395), .ZN(n10658) );
  NAND2_X2 U13905 ( .A1(aluBoi_multBoi_temppp[33]), .A2(n10659), .ZN(n12316)
         );
  XNOR2_X2 U13906 ( .A(n10660), .B(n5680), .ZN(n12213) );
  INV_X4 U13907 ( .A(n12213), .ZN(n10666) );
  NAND2_X2 U13908 ( .A1(aluBoi_multBoi_temppp[32]), .A2(n10661), .ZN(n10665)
         );
  NAND2_X2 U13909 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  NAND2_X2 U13910 ( .A1(n10665), .A2(n10664), .ZN(n12214) );
  NAND2_X2 U13911 ( .A1(n10666), .A2(n12214), .ZN(n12315) );
  XNOR2_X2 U13912 ( .A(n10667), .B(n5552), .ZN(n10668) );
  NAND2_X2 U13913 ( .A1(aluBoi_multBoi_temppp[34]), .A2(n12317), .ZN(n12318)
         );
  INV_X4 U13914 ( .A(n12318), .ZN(n10676) );
  XNOR2_X2 U13915 ( .A(n10673), .B(n10672), .ZN(n10674) );
  XNOR2_X2 U13916 ( .A(n10674), .B(n5639), .ZN(n10675) );
  OAI21_X4 U13917 ( .B1(n10677), .B2(n10676), .A(n10675), .ZN(n10870) );
  NAND2_X2 U13918 ( .A1(n10869), .A2(n10870), .ZN(n10678) );
  NAND2_X2 U13919 ( .A1(n10679), .A2(n10678), .ZN(n10680) );
  INV_X4 U13920 ( .A(n10680), .ZN(n12216) );
  NOR3_X4 U13921 ( .A1(n10681), .A2(net368481), .A3(n12216), .ZN(
        aluBoi_multBoi_N42) );
  INV_X4 U13922 ( .A(n10684), .ZN(n10685) );
  NOR2_X4 U13923 ( .A1(n10708), .A2(n10685), .ZN(n10686) );
  XNOR2_X2 U13924 ( .A(n10687), .B(n10686), .ZN(n10694) );
  INV_X4 U13925 ( .A(n10688), .ZN(n10690) );
  NAND2_X2 U13926 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NAND2_X2 U13927 ( .A1(n10692), .A2(n10691), .ZN(n10693) );
  NAND2_X2 U13928 ( .A1(n10695), .A2(net378405), .ZN(n10718) );
  NAND2_X2 U13929 ( .A1(net360904), .A2(n6541), .ZN(n10713) );
  INV_X4 U13930 ( .A(n10714), .ZN(n10843) );
  NAND4_X2 U13931 ( .A1(n10723), .A2(n9635), .A3(n10722), .A4(n10721), .ZN(
        n10771) );
  NAND2_X2 U13932 ( .A1(n10724), .A2(n10771), .ZN(n10728) );
  NOR2_X4 U13933 ( .A1(n10726), .A2(n10725), .ZN(n10727) );
  INV_X4 U13934 ( .A(n10791), .ZN(n10729) );
  NOR2_X4 U13935 ( .A1(n13706), .A2(net368209), .ZN(n10784) );
  INV_X4 U13936 ( .A(n10784), .ZN(n10730) );
  XNOR2_X2 U13937 ( .A(n10731), .B(n10730), .ZN(n10732) );
  XNOR2_X2 U13938 ( .A(n10734), .B(n10733), .ZN(n10832) );
  OAI21_X4 U13939 ( .B1(n10737), .B2(n10736), .A(n10735), .ZN(n11029) );
  NAND3_X2 U13940 ( .A1(n6435), .A2(net378405), .A3(n10738), .ZN(n10742) );
  INV_X4 U13941 ( .A(n10824), .ZN(n10739) );
  NAND3_X2 U13942 ( .A1(n10739), .A2(n6435), .A3(n10837), .ZN(n10741) );
  NAND3_X4 U13943 ( .A1(n10740), .A2(n10741), .A3(n10742), .ZN(n11030) );
  XNOR2_X2 U13944 ( .A(n10743), .B(n6541), .ZN(n10803) );
  NAND2_X2 U13945 ( .A1(net359752), .A2(n6541), .ZN(n10744) );
  OAI21_X4 U13946 ( .B1(n10803), .B2(net368185), .A(n10744), .ZN(n11028) );
  XNOR2_X2 U13947 ( .A(n10768), .B(n11028), .ZN(n10800) );
  NAND2_X2 U13948 ( .A1(net359752), .A2(n6543), .ZN(n10747) );
  XNOR2_X2 U13949 ( .A(n4997), .B(n11021), .ZN(net361537) );
  OAI22_X2 U13950 ( .A1(n10575), .A2(net368436), .B1(net368181), .B2(n10752), 
        .ZN(n10761) );
  NAND2_X2 U13951 ( .A1(n10753), .A2(n10761), .ZN(net361293) );
  NOR2_X4 U13952 ( .A1(n6001), .A2(n5761), .ZN(n10767) );
  XNOR2_X2 U13953 ( .A(n10754), .B(net361827), .ZN(n10755) );
  NAND2_X2 U13954 ( .A1(net359603), .A2(n6545), .ZN(n10758) );
  OAI21_X4 U13955 ( .B1(n10759), .B2(net368181), .A(n10758), .ZN(n10860) );
  INV_X4 U13956 ( .A(n10860), .ZN(n10764) );
  INV_X4 U13957 ( .A(n11028), .ZN(n10769) );
  NAND2_X2 U13958 ( .A1(net359752), .A2(n10724), .ZN(n10773) );
  OAI21_X4 U13959 ( .B1(net368185), .B2(n10853), .A(n10773), .ZN(net361546) );
  NAND2_X2 U13960 ( .A1(net360904), .A2(n13706), .ZN(n10777) );
  NAND2_X2 U13961 ( .A1(n10778), .A2(n10779), .ZN(n11179) );
  NAND2_X2 U13962 ( .A1(net368466), .A2(net368519), .ZN(n10787) );
  INV_X4 U13963 ( .A(n10785), .ZN(n10886) );
  INV_X4 U13964 ( .A(n10561), .ZN(n10885) );
  XNOR2_X2 U13965 ( .A(n10822), .B(n10821), .ZN(net361545) );
  XNOR2_X2 U13966 ( .A(n10795), .B(net361548), .ZN(n11031) );
  INV_X4 U13967 ( .A(n10796), .ZN(n11145) );
  NAND2_X2 U13968 ( .A1(net361825), .A2(n10855), .ZN(n10797) );
  NAND2_X2 U13969 ( .A1(n11145), .A2(n11144), .ZN(n10807) );
  NAND2_X2 U13970 ( .A1(n10801), .A2(n10807), .ZN(n10804) );
  NAND2_X2 U13971 ( .A1(net359603), .A2(n6541), .ZN(n10802) );
  OAI21_X4 U13972 ( .B1(n10803), .B2(net368181), .A(n10802), .ZN(n11147) );
  XNOR2_X2 U13973 ( .A(n10804), .B(n11147), .ZN(net361714) );
  INV_X4 U13974 ( .A(net361714), .ZN(net361291) );
  INV_X4 U13975 ( .A(n11147), .ZN(n10805) );
  INV_X4 U13976 ( .A(n10806), .ZN(n11143) );
  OAI21_X4 U13977 ( .B1(n10808), .B2(n5046), .A(n10807), .ZN(net361292) );
  NOR2_X4 U13978 ( .A1(net361808), .A2(net368462), .ZN(n10809) );
  NAND2_X2 U13979 ( .A1(net360821), .A2(n6539), .ZN(n10820) );
  NOR2_X4 U13980 ( .A1(net368209), .A2(n6539), .ZN(n10818) );
  NOR4_X2 U13981 ( .A1(n10816), .A2(n10912), .A3(n10815), .A4(n10814), .ZN(
        n10817) );
  XNOR2_X2 U13982 ( .A(n10817), .B(n10818), .ZN(n10819) );
  XNOR2_X2 U13983 ( .A(n10883), .B(n10884), .ZN(n11044) );
  NOR2_X4 U13984 ( .A1(n6387), .A2(n10985), .ZN(n10826) );
  NAND3_X4 U13985 ( .A1(n10826), .A2(n10856), .A3(n10825), .ZN(n10831) );
  NAND3_X4 U13986 ( .A1(n10831), .A2(n10991), .A3(n10830), .ZN(n11096) );
  AOI22_X2 U13987 ( .A1(n10843), .A2(n10842), .B1(n10841), .B2(n10840), .ZN(
        n10844) );
  NAND3_X4 U13988 ( .A1(n5003), .A2(n5005), .A3(n10970), .ZN(n11397) );
  NAND2_X2 U13989 ( .A1(net361524), .A2(n11095), .ZN(n10852) );
  XNOR2_X2 U13990 ( .A(n10850), .B(n10849), .ZN(n11111) );
  NAND2_X2 U13991 ( .A1(net359752), .A2(n13706), .ZN(n10851) );
  OAI21_X4 U13992 ( .B1(n11111), .B2(net368185), .A(n10851), .ZN(net361437) );
  INV_X4 U13993 ( .A(net361437), .ZN(net361756) );
  XNOR2_X2 U13994 ( .A(n10852), .B(net361756), .ZN(n11156) );
  OAI22_X2 U13995 ( .A1(n10309), .A2(net368436), .B1(net368179), .B2(n10853), 
        .ZN(n11150) );
  INV_X4 U13996 ( .A(n11150), .ZN(n10854) );
  XNOR2_X2 U13997 ( .A(n6427), .B(n10854), .ZN(n10858) );
  NAND4_X2 U13998 ( .A1(n10857), .A2(net361356), .A3(n6429), .A4(n11103), .ZN(
        n11105) );
  XNOR2_X2 U13999 ( .A(n5950), .B(n5569), .ZN(net361295) );
  XNOR2_X2 U14000 ( .A(net361740), .B(net361295), .ZN(net361312) );
  XNOR2_X2 U14001 ( .A(n10860), .B(n10859), .ZN(n10873) );
  OAI21_X4 U14002 ( .B1(n6001), .B2(n6057), .A(n10861), .ZN(n10874) );
  INV_X4 U14003 ( .A(n10863), .ZN(n10864) );
  XNOR2_X2 U14004 ( .A(n10865), .B(n10866), .ZN(n10878) );
  XNOR2_X2 U14005 ( .A(n10878), .B(n5681), .ZN(net361309) );
  NAND2_X2 U14006 ( .A1(aluBoi_multBoi_temppp[37]), .A2(n10867), .ZN(net361308) );
  AOI21_X4 U14007 ( .B1(n10870), .B2(n10869), .A(n10868), .ZN(n10877) );
  INV_X4 U14008 ( .A(n10872), .ZN(n12217) );
  XOR2_X2 U14009 ( .A(n10873), .B(aluBoi_multBoi_temppp[37]), .Z(n10875) );
  XNOR2_X2 U14010 ( .A(n10875), .B(n10874), .ZN(n12218) );
  INV_X4 U14011 ( .A(n12218), .ZN(n10876) );
  OAI21_X4 U14012 ( .B1(n10877), .B2(n12217), .A(n10876), .ZN(net361307) );
  NAND2_X2 U14013 ( .A1(net361308), .A2(net361307), .ZN(n12499) );
  NAND2_X2 U14014 ( .A1(aluBoi_multBoi_temppp[38]), .A2(n10879), .ZN(net361306) );
  INV_X4 U14015 ( .A(n10880), .ZN(n12322) );
  OAI21_X4 U14016 ( .B1(n12322), .B2(net359792), .A(net361296), .ZN(n10881) );
  OAI211_X2 U14017 ( .C1(net361709), .C2(n10881), .A(n12221), .B(net100619), 
        .ZN(n10882) );
  INV_X4 U14018 ( .A(n10882), .ZN(aluBoi_multBoi_N46) );
  NAND2_X2 U14019 ( .A1(net360821), .A2(n6537), .ZN(n10931) );
  NAND2_X2 U14020 ( .A1(n10931), .A2(n10932), .ZN(n10978) );
  XNOR2_X2 U14021 ( .A(n10887), .B(n6539), .ZN(n11116) );
  NOR2_X4 U14022 ( .A1(n10888), .A2(n10938), .ZN(n10936) );
  NOR2_X4 U14023 ( .A1(n10898), .A2(n10899), .ZN(n10900) );
  NAND3_X4 U14024 ( .A1(n10900), .A2(n10901), .A3(n10902), .ZN(n10974) );
  NAND2_X2 U14025 ( .A1(net368201), .A2(n10995), .ZN(n10908) );
  NOR2_X4 U14026 ( .A1(n10996), .A2(n10908), .ZN(n10910) );
  NAND2_X2 U14027 ( .A1(net360904), .A2(n6379), .ZN(n10973) );
  NOR3_X4 U14028 ( .A1(n10911), .A2(n10909), .A3(n10910), .ZN(n10979) );
  INV_X4 U14029 ( .A(n10917), .ZN(n10918) );
  XNOR2_X2 U14030 ( .A(n10922), .B(n10923), .ZN(n10926) );
  NAND2_X2 U14031 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  XNOR2_X2 U14032 ( .A(n10988), .B(n10987), .ZN(net361512) );
  INV_X4 U14033 ( .A(n10945), .ZN(n10935) );
  INV_X4 U14034 ( .A(n10938), .ZN(n10939) );
  AOI21_X4 U14035 ( .B1(n10944), .B2(n10943), .A(n10942), .ZN(n11118) );
  OAI22_X2 U14036 ( .A1(n9655), .A2(net368442), .B1(n5974), .B2(net368187), 
        .ZN(n10964) );
  INV_X4 U14037 ( .A(n10946), .ZN(n11117) );
  XNOR2_X2 U14038 ( .A(n10948), .B(net378128), .ZN(net361630) );
  NAND2_X2 U14039 ( .A1(n10960), .A2(n10991), .ZN(n11034) );
  INV_X4 U14040 ( .A(n10964), .ZN(n10965) );
  XNOR2_X2 U14041 ( .A(n10941), .B(n10965), .ZN(n10966) );
  XNOR2_X2 U14042 ( .A(n10967), .B(n10966), .ZN(n11124) );
  NAND2_X2 U14043 ( .A1(n11120), .A2(n11082), .ZN(n10968) );
  INV_X4 U14044 ( .A(n10968), .ZN(n11026) );
  NAND3_X4 U14045 ( .A1(n10969), .A2(n10971), .A3(n10970), .ZN(n11278) );
  INV_X4 U14046 ( .A(n10973), .ZN(n10975) );
  OAI21_X4 U14047 ( .B1(n5037), .B2(n10975), .A(n10974), .ZN(n11049) );
  NAND2_X2 U14048 ( .A1(n10978), .A2(n10977), .ZN(n10981) );
  XNOR2_X2 U14049 ( .A(n10980), .B(n10979), .ZN(n11045) );
  XNOR2_X2 U14050 ( .A(n10988), .B(n10987), .ZN(n10990) );
  OAI22_X2 U14051 ( .A1(n10995), .A2(net368446), .B1(net368187), .B2(n11102), 
        .ZN(n11011) );
  XNOR2_X2 U14052 ( .A(n10997), .B(n6535), .ZN(n11331) );
  INV_X4 U14053 ( .A(n11002), .ZN(n11070) );
  NAND2_X2 U14054 ( .A1(n11070), .A2(n11196), .ZN(n11255) );
  NAND3_X2 U14055 ( .A1(n11255), .A2(n11173), .A3(net368215), .ZN(n11006) );
  OAI21_X4 U14056 ( .B1(n5332), .B2(n11006), .A(n11005), .ZN(n11456) );
  XNOR2_X2 U14057 ( .A(n11457), .B(n11456), .ZN(n11707) );
  XNOR2_X2 U14058 ( .A(n11011), .B(n6432), .ZN(n11084) );
  INV_X4 U14059 ( .A(n11009), .ZN(n11007) );
  NAND3_X2 U14060 ( .A1(n11009), .A2(n11389), .A3(n11008), .ZN(n11017) );
  INV_X4 U14061 ( .A(n11011), .ZN(n11012) );
  NAND4_X2 U14062 ( .A1(n11018), .A2(n11017), .A3(n11016), .A4(n11015), .ZN(
        n11090) );
  INV_X4 U14063 ( .A(n11090), .ZN(n11019) );
  INV_X4 U14064 ( .A(n11021), .ZN(n11025) );
  NAND2_X2 U14065 ( .A1(n5040), .A2(n11278), .ZN(net361523) );
  NAND2_X2 U14066 ( .A1(n11155), .A2(n11130), .ZN(n11027) );
  INV_X4 U14067 ( .A(n11027), .ZN(n11113) );
  XNOR2_X2 U14068 ( .A(n11037), .B(net361443), .ZN(n11109) );
  INV_X4 U14069 ( .A(n11109), .ZN(n11152) );
  NOR2_X4 U14070 ( .A1(n5443), .A2(n5921), .ZN(n11058) );
  XNOR2_X2 U14071 ( .A(n11063), .B(n11062), .ZN(n11064) );
  NAND2_X2 U14072 ( .A1(net368201), .A2(n11173), .ZN(n11068) );
  AOI22_X2 U14073 ( .A1(n11071), .A2(n13533), .B1(n11070), .B2(n11196), .ZN(
        n11073) );
  INV_X4 U14074 ( .A(n11176), .ZN(n11072) );
  AOI21_X4 U14075 ( .B1(n11073), .B2(n11074), .A(n11072), .ZN(n11075) );
  XNOR2_X2 U14076 ( .A(n11076), .B(n11075), .ZN(n11279) );
  INV_X4 U14077 ( .A(n11082), .ZN(n11083) );
  NOR2_X4 U14078 ( .A1(n11083), .A2(net377444), .ZN(n11088) );
  INV_X4 U14079 ( .A(n11084), .ZN(n11086) );
  OAI21_X4 U14080 ( .B1(n11088), .B2(n11087), .A(n6006), .ZN(n11171) );
  INV_X4 U14081 ( .A(n11091), .ZN(n11327) );
  OAI21_X4 U14082 ( .B1(n5991), .B2(n10947), .A(n11095), .ZN(n11097) );
  OAI21_X4 U14083 ( .B1(n11098), .B2(n6071), .A(n11127), .ZN(n11099) );
  NAND3_X4 U14084 ( .A1(net376785), .A2(n11099), .A3(n11100), .ZN(net361073)
         );
  NAND2_X2 U14085 ( .A1(net359603), .A2(n6537), .ZN(n11101) );
  OAI21_X4 U14086 ( .B1(net368181), .B2(n11102), .A(n11101), .ZN(n11342) );
  XNOR2_X2 U14087 ( .A(n11343), .B(n11342), .ZN(net361008) );
  XOR2_X2 U14088 ( .A(net361008), .B(aluBoi_multBoi_temppp[44]), .Z(n11159) );
  XNOR2_X2 U14089 ( .A(n11110), .B(n11109), .ZN(net361056) );
  OAI22_X2 U14090 ( .A1(n9655), .A2(net368436), .B1(n5974), .B2(net368179), 
        .ZN(net361391) );
  OAI21_X4 U14091 ( .B1(net361400), .B2(net361401), .A(n11122), .ZN(n11119) );
  INV_X4 U14092 ( .A(net361398), .ZN(net361396) );
  OAI21_X4 U14093 ( .B1(net361396), .B2(n11120), .A(n11122), .ZN(n11121) );
  INV_X4 U14094 ( .A(n11121), .ZN(n11322) );
  NOR2_X4 U14095 ( .A1(n11323), .A2(n11322), .ZN(net361394) );
  INV_X4 U14096 ( .A(n11122), .ZN(n11123) );
  INV_X4 U14097 ( .A(net361391), .ZN(net361390) );
  NAND2_X2 U14098 ( .A1(net377443), .A2(net361386), .ZN(n11137) );
  OAI21_X4 U14099 ( .B1(n11133), .B2(n11132), .A(n11131), .ZN(n11136) );
  AOI22_X2 U14100 ( .A1(n11143), .A2(net361354), .B1(n11143), .B2(n11142), 
        .ZN(n11146) );
  XNOR2_X2 U14101 ( .A(n11148), .B(n11147), .ZN(n11149) );
  NAND2_X2 U14102 ( .A1(n5950), .A2(n11160), .ZN(n11355) );
  INV_X4 U14103 ( .A(n11355), .ZN(n11321) );
  XNOR2_X2 U14104 ( .A(n11152), .B(net361342), .ZN(n11153) );
  OAI21_X4 U14105 ( .B1(n11157), .B2(n6427), .A(n6071), .ZN(n11336) );
  XNOR2_X2 U14106 ( .A(n11337), .B(n11161), .ZN(net361318) );
  INV_X4 U14107 ( .A(net360636), .ZN(net361260) );
  AOI21_X4 U14108 ( .B1(n11162), .B2(n6009), .A(n5924), .ZN(net361275) );
  NAND2_X2 U14109 ( .A1(net361289), .A2(net361290), .ZN(n11168) );
  XNOR2_X2 U14110 ( .A(n11168), .B(n6078), .ZN(n11169) );
  NAND2_X2 U14111 ( .A1(net361260), .A2(net361261), .ZN(n11364) );
  NAND2_X2 U14112 ( .A1(n11172), .A2(n11171), .ZN(n11414) );
  NAND2_X2 U14113 ( .A1(n11255), .A2(n11173), .ZN(n11177) );
  INV_X4 U14114 ( .A(n11177), .ZN(n11174) );
  NAND2_X2 U14115 ( .A1(n11174), .A2(n5983), .ZN(n11263) );
  OAI22_X2 U14116 ( .A1(n11067), .A2(net368447), .B1(net368187), .B2(n11263), 
        .ZN(n11417) );
  INV_X4 U14117 ( .A(n11208), .ZN(n11178) );
  AOI21_X4 U14118 ( .B1(n11176), .B2(net368195), .A(n11076), .ZN(n11214) );
  NOR2_X4 U14119 ( .A1(n11178), .A2(n11207), .ZN(n11203) );
  NAND2_X2 U14120 ( .A1(net360821), .A2(n6529), .ZN(n11219) );
  INV_X4 U14121 ( .A(n11185), .ZN(n11237) );
  NAND2_X2 U14122 ( .A1(net368201), .A2(n11199), .ZN(n11200) );
  XNOR2_X2 U14123 ( .A(n11226), .B(n11225), .ZN(n11216) );
  INV_X4 U14124 ( .A(n11216), .ZN(n11202) );
  XNOR2_X2 U14125 ( .A(n11203), .B(n11202), .ZN(n11416) );
  XNOR2_X2 U14126 ( .A(n11417), .B(n11216), .ZN(n11211) );
  XNOR2_X2 U14127 ( .A(n11211), .B(n11210), .ZN(n11418) );
  NAND3_X4 U14128 ( .A1(net361073), .A2(n11409), .A3(n11327), .ZN(n11258) );
  OAI21_X4 U14129 ( .B1(n5923), .B2(n11212), .A(n6164), .ZN(n11333) );
  NAND2_X2 U14130 ( .A1(n11311), .A2(n6529), .ZN(n11234) );
  INV_X4 U14131 ( .A(n11233), .ZN(n11527) );
  NAND2_X2 U14132 ( .A1(n11527), .A2(n11298), .ZN(n11312) );
  INV_X4 U14133 ( .A(n11238), .ZN(n11240) );
  NAND2_X2 U14134 ( .A1(net360904), .A2(n6529), .ZN(n11239) );
  OAI21_X4 U14135 ( .B1(n11241), .B2(n11240), .A(n11239), .ZN(n11371) );
  INV_X4 U14136 ( .A(n11371), .ZN(n11471) );
  NAND2_X2 U14137 ( .A1(net360821), .A2(n6527), .ZN(n11284) );
  INV_X4 U14138 ( .A(n11284), .ZN(n11252) );
  INV_X4 U14139 ( .A(n11246), .ZN(n11292) );
  NAND2_X2 U14140 ( .A1(n11284), .A2(net368211), .ZN(n11251) );
  OAI21_X4 U14141 ( .B1(n6058), .B2(n11252), .A(n11251), .ZN(n11470) );
  XNOR2_X2 U14142 ( .A(n11471), .B(n11253), .ZN(n11643) );
  OAI22_X2 U14143 ( .A1(n11256), .A2(net368444), .B1(n11315), .B2(net368187), 
        .ZN(n11274) );
  INV_X4 U14144 ( .A(n11418), .ZN(n11736) );
  NAND2_X2 U14145 ( .A1(n11261), .A2(n11335), .ZN(net361027) );
  OAI21_X4 U14146 ( .B1(net368181), .B2(n11263), .A(n11262), .ZN(net361028) );
  NOR2_X4 U14147 ( .A1(n11265), .A2(n11266), .ZN(n11272) );
  INV_X4 U14148 ( .A(n11269), .ZN(n11270) );
  INV_X4 U14149 ( .A(n11277), .ZN(n11290) );
  OAI21_X4 U14150 ( .B1(n11394), .B2(n11281), .A(n11280), .ZN(n11289) );
  NAND2_X2 U14151 ( .A1(n6423), .A2(n11282), .ZN(n11391) );
  INV_X4 U14152 ( .A(n11391), .ZN(n11287) );
  INV_X4 U14153 ( .A(n5034), .ZN(n11285) );
  AOI21_X4 U14154 ( .B1(n11287), .B2(n11286), .A(n11285), .ZN(n11288) );
  OAI21_X4 U14155 ( .B1(n11290), .B2(n11289), .A(n11288), .ZN(n11426) );
  NAND2_X2 U14156 ( .A1(n11292), .A2(n11291), .ZN(n11293) );
  NAND2_X2 U14157 ( .A1(net360904), .A2(n6527), .ZN(n11294) );
  OAI21_X4 U14158 ( .B1(n11295), .B2(net368195), .A(n11294), .ZN(n11386) );
  NAND2_X2 U14159 ( .A1(net360821), .A2(n6525), .ZN(n11309) );
  NAND3_X2 U14160 ( .A1(n11378), .A2(n11483), .A3(net368215), .ZN(n11308) );
  XNOR2_X2 U14161 ( .A(n11386), .B(n11385), .ZN(n11425) );
  OAI22_X2 U14162 ( .A1(n11191), .A2(net368446), .B1(net368187), .B2(n11431), 
        .ZN(n11427) );
  OAI22_X2 U14163 ( .A1(n11316), .A2(net368436), .B1(n11315), .B2(net368179), 
        .ZN(n11433) );
  INV_X4 U14164 ( .A(n11433), .ZN(n11317) );
  AOI21_X4 U14165 ( .B1(n11321), .B2(n11354), .A(n11358), .ZN(n11326) );
  NOR2_X4 U14166 ( .A1(n11323), .A2(n11322), .ZN(net361083) );
  INV_X4 U14167 ( .A(n11357), .ZN(n11325) );
  NOR2_X4 U14168 ( .A1(n11326), .A2(n11325), .ZN(n11351) );
  NAND3_X4 U14169 ( .A1(n11261), .A2(n11335), .A3(net361028), .ZN(net361031)
         );
  INV_X4 U14170 ( .A(n11342), .ZN(n11344) );
  NAND2_X2 U14171 ( .A1(n11344), .A2(n11343), .ZN(n11352) );
  NAND3_X4 U14172 ( .A1(n11348), .A2(net361022), .A3(net361031), .ZN(n11349)
         );
  OAI21_X4 U14173 ( .B1(n11351), .B2(n11350), .A(n11349), .ZN(net360927) );
  INV_X4 U14174 ( .A(net361020), .ZN(net361033) );
  XNOR2_X2 U14175 ( .A(net361027), .B(net361028), .ZN(net361019) );
  INV_X4 U14176 ( .A(n12327), .ZN(n11370) );
  XNOR2_X2 U14177 ( .A(net361018), .B(net361019), .ZN(n11368) );
  XNOR2_X2 U14178 ( .A(n11368), .B(n5646), .ZN(n11360) );
  XNOR2_X2 U14179 ( .A(n11362), .B(net361008), .ZN(n11363) );
  INV_X4 U14180 ( .A(net361009), .ZN(net359918) );
  XNOR2_X2 U14181 ( .A(net378491), .B(n5560), .ZN(net359919) );
  NAND2_X2 U14182 ( .A1(n11471), .A2(n11470), .ZN(n11465) );
  NAND3_X4 U14183 ( .A1(n11374), .A2(n5939), .A3(n11373), .ZN(n11594) );
  NAND3_X4 U14184 ( .A1(n11627), .A2(n5202), .A3(n11465), .ZN(n11458) );
  INV_X4 U14185 ( .A(n6525), .ZN(n11379) );
  NAND2_X2 U14186 ( .A1(net360821), .A2(n6523), .ZN(n11443) );
  INV_X4 U14187 ( .A(n11443), .ZN(n11381) );
  AOI21_X4 U14188 ( .B1(net368215), .B2(n11382), .A(n11381), .ZN(n11383) );
  XNOR2_X2 U14189 ( .A(n11384), .B(n11383), .ZN(n11467) );
  XNOR2_X2 U14190 ( .A(n11407), .B(n11440), .ZN(n11700) );
  INV_X4 U14191 ( .A(n11408), .ZN(n11413) );
  NAND2_X2 U14192 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  NAND2_X2 U14193 ( .A1(n11415), .A2(n11414), .ZN(n11423) );
  INV_X4 U14194 ( .A(n11419), .ZN(n11493) );
  XNOR2_X2 U14195 ( .A(n11426), .B(n6106), .ZN(n11428) );
  NAND2_X2 U14196 ( .A1(n11513), .A2(n11512), .ZN(n11508) );
  NAND2_X2 U14197 ( .A1(net359603), .A2(n6529), .ZN(n11430) );
  OAI21_X4 U14198 ( .B1(net368181), .B2(n11431), .A(n11430), .ZN(n11516) );
  XNOR2_X2 U14199 ( .A(n11515), .B(n11516), .ZN(n11674) );
  XNOR2_X2 U14200 ( .A(n11436), .B(n5141), .ZN(n11669) );
  OAI21_X4 U14201 ( .B1(net360915), .B2(n12328), .A(n11437), .ZN(net359915) );
  AOI211_X4 U14202 ( .C1(n11438), .C2(n6069), .A(net368481), .B(net360914), 
        .ZN(aluBoi_multBoi_N54) );
  INV_X4 U14203 ( .A(n11439), .ZN(n11442) );
  NAND2_X2 U14204 ( .A1(n11495), .A2(n11738), .ZN(n11491) );
  NAND2_X2 U14205 ( .A1(n11443), .A2(net368211), .ZN(n11446) );
  NAND2_X2 U14206 ( .A1(n6083), .A2(n11443), .ZN(n11444) );
  NAND2_X2 U14207 ( .A1(net360904), .A2(n6523), .ZN(n11461) );
  NAND2_X2 U14208 ( .A1(net360821), .A2(n6521), .ZN(n11448) );
  INV_X4 U14209 ( .A(n11502), .ZN(n11449) );
  XNOR2_X2 U14210 ( .A(n6552), .B(n11449), .ZN(n11702) );
  XNOR2_X2 U14211 ( .A(n11450), .B(n6092), .ZN(n11688) );
  INV_X4 U14212 ( .A(n11688), .ZN(n11452) );
  NAND2_X2 U14213 ( .A1(net359603), .A2(n6527), .ZN(n11451) );
  INV_X4 U14214 ( .A(n6525), .ZN(n11454) );
  INV_X4 U14215 ( .A(n11641), .ZN(n11455) );
  NAND2_X2 U14216 ( .A1(n6108), .A2(n5893), .ZN(n11573) );
  NOR2_X4 U14217 ( .A1(n11467), .A2(n11464), .ZN(n11466) );
  NAND2_X2 U14218 ( .A1(n11471), .A2(n5998), .ZN(n11595) );
  INV_X4 U14219 ( .A(n11595), .ZN(n11472) );
  OAI21_X4 U14220 ( .B1(n11474), .B2(n11644), .A(n11473), .ZN(n11551) );
  INV_X4 U14221 ( .A(n11551), .ZN(n11534) );
  OAI21_X4 U14222 ( .B1(n6553), .B2(n11475), .A(n5893), .ZN(n11572) );
  INV_X4 U14223 ( .A(n11607), .ZN(n11479) );
  NAND2_X2 U14224 ( .A1(net360821), .A2(n6519), .ZN(n11481) );
  OAI21_X4 U14225 ( .B1(n11482), .B2(net368209), .A(n11481), .ZN(n11536) );
  INV_X4 U14226 ( .A(n11536), .ZN(n11588) );
  NAND2_X2 U14227 ( .A1(n6063), .A2(n6521), .ZN(n11485) );
  OAI21_X4 U14228 ( .B1(n11487), .B2(net368462), .A(n11486), .ZN(n11537) );
  INV_X4 U14229 ( .A(n11537), .ZN(n11587) );
  XNOR2_X2 U14230 ( .A(n11588), .B(n11587), .ZN(n11582) );
  INV_X4 U14231 ( .A(n6523), .ZN(n11488) );
  OAI22_X2 U14232 ( .A1(n11488), .A2(net368446), .B1(n6083), .B2(net368187), 
        .ZN(n11558) );
  XNOR2_X2 U14233 ( .A(n11582), .B(n11558), .ZN(n11574) );
  XNOR2_X2 U14234 ( .A(n11489), .B(n11574), .ZN(n11506) );
  NOR3_X4 U14235 ( .A1(n11742), .A2(n11741), .A3(n11496), .ZN(n11497) );
  XNOR2_X2 U14236 ( .A(n11501), .B(n6553), .ZN(n11503) );
  INV_X4 U14237 ( .A(n11506), .ZN(n11560) );
  INV_X4 U14238 ( .A(n11516), .ZN(n11510) );
  OAI21_X4 U14239 ( .B1(n11511), .B2(n6128), .A(n11510), .ZN(n11912) );
  INV_X4 U14240 ( .A(n11515), .ZN(n11517) );
  NAND2_X2 U14241 ( .A1(net360821), .A2(net368572), .ZN(n11526) );
  NAND2_X2 U14242 ( .A1(n11522), .A2(net368572), .ZN(n11606) );
  NAND3_X2 U14243 ( .A1(n11605), .A2(n11606), .A3(net368215), .ZN(n11525) );
  NAND2_X2 U14244 ( .A1(n11526), .A2(n11525), .ZN(n11619) );
  INV_X4 U14245 ( .A(n11619), .ZN(n11616) );
  XNOR2_X2 U14246 ( .A(n11616), .B(n11615), .ZN(n11637) );
  INV_X4 U14247 ( .A(n11637), .ZN(n11589) );
  INV_X4 U14248 ( .A(n6521), .ZN(n11532) );
  OAI22_X2 U14249 ( .A1(n11532), .A2(net368447), .B1(net368187), .B2(n11655), 
        .ZN(n11584) );
  INV_X4 U14250 ( .A(n11584), .ZN(n11751) );
  NOR2_X4 U14251 ( .A1(n6553), .A2(n11556), .ZN(n11535) );
  INV_X4 U14252 ( .A(n11535), .ZN(n11540) );
  NAND2_X2 U14253 ( .A1(n11582), .A2(n11614), .ZN(n11542) );
  AOI21_X4 U14254 ( .B1(n11541), .B2(n11540), .A(n11539), .ZN(n11570) );
  INV_X4 U14255 ( .A(n11542), .ZN(n11543) );
  NAND2_X2 U14256 ( .A1(net359603), .A2(n6523), .ZN(n11545) );
  OAI21_X4 U14257 ( .B1(n6083), .B2(net368179), .A(n11545), .ZN(n11892) );
  INV_X4 U14258 ( .A(n11613), .ZN(n11552) );
  OAI21_X4 U14259 ( .B1(n6553), .B2(n11556), .A(n11555), .ZN(n11579) );
  XNOR2_X2 U14260 ( .A(n11561), .B(n11562), .ZN(n12121) );
  INV_X4 U14261 ( .A(n11565), .ZN(n11684) );
  INV_X4 U14262 ( .A(n11960), .ZN(n12119) );
  XNOR2_X2 U14263 ( .A(n5186), .B(n11561), .ZN(n11893) );
  XNOR2_X2 U14264 ( .A(n11544), .B(n11571), .ZN(n11701) );
  XNOR2_X2 U14265 ( .A(n11575), .B(n11574), .ZN(n11576) );
  NAND2_X2 U14266 ( .A1(n11869), .A2(n11870), .ZN(n11897) );
  OAI21_X4 U14267 ( .B1(n11863), .B2(net368185), .A(n11585), .ZN(n11760) );
  INV_X4 U14268 ( .A(n11760), .ZN(n11848) );
  NAND2_X2 U14269 ( .A1(n11588), .A2(n11587), .ZN(n11639) );
  AOI21_X4 U14270 ( .B1(n11713), .B2(n11602), .A(n6553), .ZN(n11604) );
  INV_X4 U14271 ( .A(net368572), .ZN(net360723) );
  NAND2_X2 U14272 ( .A1(n11614), .A2(n11613), .ZN(n11618) );
  OAI21_X4 U14273 ( .B1(n11622), .B2(n11827), .A(n11621), .ZN(n11752) );
  INV_X4 U14274 ( .A(n11628), .ZN(n11630) );
  AOI21_X4 U14275 ( .B1(n11798), .B2(n11648), .A(n11824), .ZN(n11649) );
  OAI21_X4 U14276 ( .B1(n11651), .B2(n11650), .A(n11649), .ZN(n11714) );
  NAND2_X2 U14277 ( .A1(net359603), .A2(n6521), .ZN(n11654) );
  OAI21_X4 U14278 ( .B1(net368181), .B2(n11655), .A(n11654), .ZN(n11914) );
  INV_X4 U14279 ( .A(n11914), .ZN(n11656) );
  XNOR2_X2 U14280 ( .A(n5880), .B(n11656), .ZN(n11663) );
  INV_X4 U14281 ( .A(n11849), .ZN(n11858) );
  NOR4_X2 U14282 ( .A1(n6207), .A2(n11660), .A3(n11659), .A4(n6092), .ZN(
        n11661) );
  INV_X4 U14283 ( .A(n11897), .ZN(n11662) );
  XNOR2_X2 U14284 ( .A(n6082), .B(n11687), .ZN(n11686) );
  INV_X4 U14285 ( .A(n11665), .ZN(n11680) );
  XNOR2_X2 U14286 ( .A(n11666), .B(n11684), .ZN(n11679) );
  XNOR2_X2 U14287 ( .A(n11679), .B(aluBoi_multBoi_temppp[50]), .ZN(n11667) );
  INV_X4 U14288 ( .A(n12508), .ZN(n12506) );
  NAND2_X2 U14289 ( .A1(n5560), .A2(net378491), .ZN(n11670) );
  NAND3_X2 U14290 ( .A1(net360639), .A2(n11671), .A3(net359916), .ZN(n11672)
         );
  INV_X4 U14291 ( .A(n11674), .ZN(n11678) );
  XNOR2_X2 U14292 ( .A(n11680), .B(n11679), .ZN(n11681) );
  INV_X4 U14293 ( .A(n11687), .ZN(n11689) );
  INV_X4 U14294 ( .A(n12121), .ZN(n11955) );
  INV_X4 U14295 ( .A(n11698), .ZN(aluBoi_multBoi_N58) );
  AOI21_X4 U14296 ( .B1(n11512), .B2(n11738), .A(n11701), .ZN(n11705) );
  INV_X4 U14297 ( .A(n5309), .ZN(n11731) );
  NAND4_X2 U14298 ( .A1(n6374), .A2(net360550), .A3(n11729), .A4(n11728), .ZN(
        n11724) );
  XNOR2_X2 U14299 ( .A(n11775), .B(n5895), .ZN(n11778) );
  INV_X4 U14300 ( .A(n5996), .ZN(n11748) );
  NOR2_X4 U14301 ( .A1(n11741), .A2(n11735), .ZN(n11739) );
  NAND3_X4 U14302 ( .A1(n11737), .A2(n11738), .A3(n11739), .ZN(n11747) );
  OAI21_X4 U14303 ( .B1(n11745), .B2(n11744), .A(n11743), .ZN(n11746) );
  NAND3_X4 U14304 ( .A1(n11748), .A2(n11747), .A3(n11746), .ZN(n11749) );
  NOR2_X4 U14305 ( .A1(n11756), .A2(n11757), .ZN(n11759) );
  INV_X4 U14306 ( .A(n6517), .ZN(n11764) );
  XNOR2_X2 U14307 ( .A(n11765), .B(n6517), .ZN(n12020) );
  NOR2_X4 U14308 ( .A1(n11767), .A2(net329432), .ZN(n11773) );
  XNOR2_X2 U14309 ( .A(n11813), .B(n11814), .ZN(n11822) );
  INV_X4 U14310 ( .A(n11822), .ZN(n11808) );
  XNOR2_X2 U14311 ( .A(n11808), .B(n11790), .ZN(n11782) );
  INV_X4 U14312 ( .A(n5309), .ZN(n11776) );
  XNOR2_X2 U14313 ( .A(n5890), .B(n11780), .ZN(n11785) );
  XNOR2_X2 U14314 ( .A(n11782), .B(n11781), .ZN(n11999) );
  NAND2_X2 U14315 ( .A1(n11999), .A2(n5919), .ZN(n12012) );
  XNOR2_X2 U14316 ( .A(n11788), .B(n5894), .ZN(n11784) );
  XNOR2_X2 U14317 ( .A(n11789), .B(n11808), .ZN(n11791) );
  NOR2_X4 U14318 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  OAI21_X4 U14319 ( .B1(n11795), .B2(n12012), .A(n11794), .ZN(n12004) );
  INV_X4 U14320 ( .A(n12004), .ZN(n12194) );
  NAND2_X2 U14321 ( .A1(n11806), .A2(n11796), .ZN(n11817) );
  INV_X4 U14322 ( .A(n11817), .ZN(n11804) );
  INV_X4 U14323 ( .A(n11805), .ZN(n11807) );
  OAI22_X2 U14324 ( .A1(net360445), .A2(net368462), .B1(net360206), .B2(
        net368195), .ZN(n11984) );
  XNOR2_X2 U14325 ( .A(n6027), .B(n6515), .ZN(n12064) );
  XNOR2_X2 U14326 ( .A(n11984), .B(n11983), .ZN(n12040) );
  NAND2_X2 U14327 ( .A1(n12040), .A2(n11820), .ZN(n11830) );
  OAI21_X4 U14328 ( .B1(n11822), .B2(n11821), .A(n11820), .ZN(n11823) );
  NOR3_X4 U14329 ( .A1(n12041), .A2(n12040), .A3(n12043), .ZN(n11829) );
  NOR2_X4 U14330 ( .A1(n6385), .A2(n11824), .ZN(n11826) );
  INV_X4 U14331 ( .A(n12011), .ZN(n11987) );
  INV_X4 U14332 ( .A(n11986), .ZN(n12010) );
  XNOR2_X2 U14333 ( .A(n11987), .B(n12010), .ZN(n12190) );
  NAND2_X2 U14334 ( .A1(net359603), .A2(n5309), .ZN(n11832) );
  NAND2_X2 U14335 ( .A1(net359603), .A2(net368572), .ZN(n11846) );
  OAI21_X4 U14336 ( .B1(net368181), .B2(net360403), .A(n11846), .ZN(n11928) );
  NAND3_X4 U14337 ( .A1(n11884), .A2(n11928), .A3(n11885), .ZN(n12112) );
  NAND2_X2 U14338 ( .A1(n11850), .A2(n11855), .ZN(n11851) );
  OAI22_X2 U14339 ( .A1(n5305), .A2(net368436), .B1(n11863), .B2(net368179), 
        .ZN(n11900) );
  XNOR2_X2 U14340 ( .A(n11864), .B(n5995), .ZN(n11899) );
  NAND2_X2 U14341 ( .A1(n11900), .A2(n11899), .ZN(n11944) );
  NAND2_X2 U14342 ( .A1(n11997), .A2(n11998), .ZN(n11889) );
  INV_X4 U14343 ( .A(n6430), .ZN(n11883) );
  OAI22_X2 U14344 ( .A1(net360360), .A2(net368436), .B1(n4987), .B2(net368179), 
        .ZN(n11890) );
  INV_X4 U14345 ( .A(n11890), .ZN(n11882) );
  XNOR2_X2 U14346 ( .A(n11903), .B(n5403), .ZN(n12095) );
  INV_X4 U14347 ( .A(n11929), .ZN(n11886) );
  NOR3_X4 U14348 ( .A1(n11888), .A2(n12095), .A3(n11887), .ZN(n12087) );
  NAND4_X2 U14349 ( .A1(n11901), .A2(n11907), .A3(n12112), .A4(n11902), .ZN(
        n11906) );
  NAND4_X2 U14350 ( .A1(n11907), .A2(n12120), .A3(n12112), .A4(n11902), .ZN(
        n11905) );
  XNOR2_X2 U14351 ( .A(n11903), .B(n5403), .ZN(n12118) );
  INV_X4 U14352 ( .A(n11928), .ZN(n11908) );
  NAND2_X2 U14353 ( .A1(n11908), .A2(n11929), .ZN(n11909) );
  OAI21_X4 U14354 ( .B1(n11910), .B2(n5884), .A(n11909), .ZN(n12113) );
  XNOR2_X2 U14355 ( .A(n12145), .B(n12146), .ZN(net359520) );
  INV_X4 U14356 ( .A(n11912), .ZN(n11918) );
  NAND2_X2 U14357 ( .A1(n11901), .A2(n11945), .ZN(n11921) );
  NAND2_X2 U14358 ( .A1(n11960), .A2(n11955), .ZN(n11932) );
  XNOR2_X2 U14359 ( .A(n11929), .B(n11928), .ZN(n11947) );
  XNOR2_X2 U14360 ( .A(n11930), .B(n6013), .ZN(net360254) );
  INV_X4 U14361 ( .A(n11932), .ZN(n11934) );
  XNOR2_X2 U14362 ( .A(n11937), .B(n5551), .ZN(net360265) );
  XNOR2_X2 U14363 ( .A(n11939), .B(n11938), .ZN(net360262) );
  NAND2_X2 U14364 ( .A1(net360261), .A2(net360262), .ZN(net359532) );
  INV_X4 U14365 ( .A(n12519), .ZN(n11970) );
  INV_X4 U14366 ( .A(n11946), .ZN(n11952) );
  INV_X4 U14367 ( .A(n11954), .ZN(n12033) );
  INV_X4 U14368 ( .A(n11962), .ZN(n11966) );
  OAI21_X4 U14369 ( .B1(n11966), .B2(n11965), .A(n11964), .ZN(n11967) );
  NAND2_X2 U14370 ( .A1(n11967), .A2(n11969), .ZN(n12147) );
  XNOR2_X2 U14371 ( .A(n12149), .B(n5537), .ZN(n12332) );
  INV_X4 U14372 ( .A(net359678), .ZN(n12518) );
  INV_X4 U14373 ( .A(n11972), .ZN(n12335) );
  NOR3_X4 U14374 ( .A1(n11973), .A2(net368481), .A3(n12335), .ZN(
        aluBoi_multBoi_N62) );
  OAI21_X4 U14375 ( .B1(net368181), .B2(net360206), .A(n11974), .ZN(n12105) );
  INV_X4 U14376 ( .A(n6515), .ZN(n11975) );
  INV_X4 U14377 ( .A(n6513), .ZN(n11982) );
  OAI21_X4 U14378 ( .B1(n11980), .B2(n11979), .A(n6513), .ZN(n11981) );
  XNOR2_X2 U14379 ( .A(n5966), .B(n11995), .ZN(n12042) );
  NAND2_X2 U14380 ( .A1(n11985), .A2(net360198), .ZN(n12074) );
  NAND2_X2 U14381 ( .A1(n5042), .A2(n11988), .ZN(n12022) );
  INV_X4 U14382 ( .A(net360198), .ZN(net360197) );
  XNOR2_X2 U14383 ( .A(n11996), .B(net360197), .ZN(n11990) );
  NAND2_X2 U14384 ( .A1(n6428), .A2(n12074), .ZN(n12005) );
  INV_X4 U14385 ( .A(n6513), .ZN(n11991) );
  INV_X4 U14386 ( .A(n6511), .ZN(n11993) );
  XNOR2_X2 U14387 ( .A(n12047), .B(n12048), .ZN(n12071) );
  INV_X4 U14388 ( .A(n12071), .ZN(n12172) );
  NAND2_X2 U14389 ( .A1(net359752), .A2(n6515), .ZN(n11994) );
  INV_X4 U14390 ( .A(n12273), .ZN(n12162) );
  OAI21_X4 U14391 ( .B1(n6097), .B2(n11996), .A(n12167), .ZN(n12067) );
  XNOR2_X2 U14392 ( .A(n12067), .B(n12068), .ZN(n12165) );
  INV_X4 U14393 ( .A(n12021), .ZN(n12002) );
  NAND2_X2 U14394 ( .A1(n6430), .A2(n11998), .ZN(n12000) );
  INV_X4 U14395 ( .A(n12074), .ZN(n12003) );
  OAI21_X4 U14396 ( .B1(n12008), .B2(n12007), .A(n12006), .ZN(n12104) );
  NAND2_X2 U14397 ( .A1(n12011), .A2(n12010), .ZN(n12017) );
  INV_X4 U14398 ( .A(n12012), .ZN(n12013) );
  NAND2_X2 U14399 ( .A1(n12015), .A2(n12016), .ZN(n12025) );
  NAND2_X2 U14400 ( .A1(n12017), .A2(n12025), .ZN(n12199) );
  XNOR2_X2 U14401 ( .A(n12018), .B(n6399), .ZN(n12115) );
  NAND2_X2 U14402 ( .A1(net359603), .A2(n6517), .ZN(n12019) );
  OAI21_X4 U14403 ( .B1(n12246), .B2(n12245), .A(n12244), .ZN(n12423) );
  NAND2_X2 U14404 ( .A1(n12190), .A2(n12025), .ZN(n12434) );
  NAND3_X4 U14405 ( .A1(n12434), .A2(n12435), .A3(n5266), .ZN(n12465) );
  INV_X4 U14406 ( .A(n12465), .ZN(n12027) );
  XNOR2_X2 U14407 ( .A(n12027), .B(n12026), .ZN(n12109) );
  INV_X4 U14408 ( .A(n12109), .ZN(n12085) );
  NOR2_X4 U14409 ( .A1(n12032), .A2(n12094), .ZN(n12034) );
  OAI21_X4 U14410 ( .B1(n12037), .B2(n12036), .A(n12035), .ZN(n12419) );
  OAI22_X2 U14411 ( .A1(n11991), .A2(net368444), .B1(net368187), .B2(n12204), 
        .ZN(n12163) );
  INV_X4 U14412 ( .A(n12163), .ZN(n12052) );
  INV_X4 U14413 ( .A(n12175), .ZN(n12062) );
  INV_X4 U14414 ( .A(n12176), .ZN(n12061) );
  XNOR2_X2 U14415 ( .A(n12062), .B(n12061), .ZN(n12349) );
  XNOR2_X2 U14416 ( .A(n12063), .B(n5971), .ZN(n12271) );
  INV_X4 U14417 ( .A(n12157), .ZN(n12065) );
  XNOR2_X2 U14418 ( .A(n12358), .B(n12065), .ZN(n12066) );
  INV_X4 U14419 ( .A(n12066), .ZN(n12239) );
  XNOR2_X2 U14420 ( .A(n12067), .B(n12068), .ZN(n12270) );
  XNOR2_X2 U14421 ( .A(n12072), .B(n5914), .ZN(n12161) );
  INV_X4 U14422 ( .A(n12161), .ZN(n12275) );
  INV_X4 U14423 ( .A(n12076), .ZN(n12077) );
  NOR2_X4 U14424 ( .A1(n12077), .A2(n12078), .ZN(n12080) );
  XNOR2_X2 U14425 ( .A(n12238), .B(n12239), .ZN(n12406) );
  XNOR2_X2 U14426 ( .A(aluBoi_multBoi_temppp[59]), .B(n12304), .ZN(n12082) );
  XNOR2_X2 U14427 ( .A(n12083), .B(n12082), .ZN(n12336) );
  XNOR2_X2 U14428 ( .A(n12404), .B(n12304), .ZN(n12084) );
  NAND2_X2 U14429 ( .A1(n12532), .A2(net359501), .ZN(n12152) );
  NAND2_X2 U14430 ( .A1(n12092), .A2(n12133), .ZN(n12151) );
  NAND2_X2 U14431 ( .A1(n6155), .A2(n11834), .ZN(n12110) );
  XNOR2_X2 U14432 ( .A(n12106), .B(n12105), .ZN(n12285) );
  OAI21_X4 U14433 ( .B1(n12292), .B2(n6431), .A(n12107), .ZN(n12289) );
  NAND2_X2 U14434 ( .A1(n12290), .A2(n5134), .ZN(n12141) );
  INV_X4 U14435 ( .A(n12110), .ZN(n12111) );
  INV_X4 U14436 ( .A(n12114), .ZN(n12117) );
  NAND4_X2 U14437 ( .A1(n12122), .A2(n12125), .A3(n12123), .A4(n12124), .ZN(
        n12126) );
  INV_X4 U14438 ( .A(n12126), .ZN(n12294) );
  XNOR2_X2 U14439 ( .A(n12131), .B(n12285), .ZN(net360017) );
  INV_X4 U14440 ( .A(aluBoi_multBoi_temppp[58]), .ZN(n12144) );
  NAND2_X2 U14441 ( .A1(n12132), .A2(n12144), .ZN(n12530) );
  XNOR2_X2 U14442 ( .A(n12145), .B(n12291), .ZN(n12139) );
  XNOR2_X2 U14443 ( .A(n12149), .B(n5537), .ZN(net359678) );
  INV_X4 U14444 ( .A(n12244), .ZN(n12287) );
  OAI211_X2 U14445 ( .C1(n12287), .C2(n12285), .A(n12406), .B(n12159), .ZN(
        n12377) );
  INV_X4 U14446 ( .A(n12349), .ZN(n12256) );
  INV_X4 U14447 ( .A(n6511), .ZN(n12166) );
  INV_X4 U14448 ( .A(n12168), .ZN(n12169) );
  NAND2_X2 U14449 ( .A1(n12176), .A2(n12175), .ZN(n12259) );
  INV_X4 U14450 ( .A(n12259), .ZN(n12177) );
  OAI21_X4 U14451 ( .B1(n12181), .B2(n12180), .A(n12179), .ZN(n12263) );
  INV_X4 U14452 ( .A(n12263), .ZN(n12188) );
  OAI22_X2 U14453 ( .A1(n12185), .A2(net368462), .B1(net368195), .B2(n12342), 
        .ZN(n12250) );
  INV_X4 U14454 ( .A(n12250), .ZN(n12186) );
  XNOR2_X2 U14455 ( .A(n12187), .B(n12186), .ZN(n12254) );
  INV_X4 U14456 ( .A(n12254), .ZN(n12264) );
  OAI211_X2 U14457 ( .C1(n12196), .C2(n12195), .A(n12369), .B(n5957), .ZN(
        n12232) );
  NAND2_X2 U14458 ( .A1(net359603), .A2(n6513), .ZN(n12203) );
  XNOR2_X2 U14459 ( .A(n12301), .B(net359418), .ZN(n12536) );
  XNOR2_X2 U14460 ( .A(n12537), .B(n12536), .ZN(n12528) );
  MUX2_X2 U14461 ( .A(aluBoi_multBoi_temppp[26]), .B(n12207), .S(net367631), 
        .Z(n13678) );
  MUX2_X2 U14462 ( .A(aluBoi_multBoi_temppp[25]), .B(n12208), .S(net367631), 
        .Z(n13681) );
  MUX2_X2 U14463 ( .A(n12212), .B(n12211), .S(net367631), .Z(
        aluBoi_multBoi_N35) );
  XNOR2_X2 U14464 ( .A(n12214), .B(n12213), .ZN(n12215) );
  NOR2_X4 U14465 ( .A1(n12217), .A2(n12216), .ZN(n12219) );
  XNOR2_X2 U14466 ( .A(n12219), .B(n12218), .ZN(n12220) );
  NOR2_X4 U14467 ( .A1(net367631), .A2(n12220), .ZN(aluBoi_multBoi_N43) );
  XNOR2_X2 U14468 ( .A(n12324), .B(net375948), .ZN(n12222) );
  XNOR2_X2 U14469 ( .A(net359918), .B(net359919), .ZN(n12223) );
  NAND2_X2 U14470 ( .A1(aluBoi_multBoi_temppp[52]), .A2(net359911), .ZN(n12509) );
  XNOR2_X2 U14471 ( .A(n12226), .B(net377454), .ZN(n12227) );
  NOR2_X4 U14472 ( .A1(net368481), .A2(n12227), .ZN(aluBoi_multBoi_N59) );
  NOR2_X4 U14473 ( .A1(n12518), .A2(n5048), .ZN(n12229) );
  INV_X4 U14474 ( .A(net359905), .ZN(net359515) );
  XNOR2_X2 U14475 ( .A(n12230), .B(net359765), .ZN(n12231) );
  NOR2_X4 U14476 ( .A1(n12234), .A2(n12408), .ZN(n12235) );
  INV_X4 U14477 ( .A(n6511), .ZN(n12249) );
  OAI22_X2 U14478 ( .A1(n12249), .A2(net368436), .B1(n6049), .B2(net368179), 
        .ZN(n12382) );
  INV_X4 U14479 ( .A(n12354), .ZN(n12344) );
  INV_X4 U14480 ( .A(n12460), .ZN(n12568) );
  NAND2_X2 U14481 ( .A1(n12254), .A2(n12354), .ZN(n12257) );
  NAND2_X2 U14482 ( .A1(n12568), .A2(n12257), .ZN(n12258) );
  INV_X4 U14483 ( .A(n12258), .ZN(n12350) );
  NAND2_X2 U14484 ( .A1(n12354), .A2(n12259), .ZN(n12351) );
  NAND2_X2 U14485 ( .A1(n12350), .A2(n12351), .ZN(n12261) );
  NAND2_X2 U14486 ( .A1(n12344), .A2(n12265), .ZN(n12268) );
  OAI21_X4 U14487 ( .B1(net368185), .B2(n12342), .A(n12269), .ZN(n12427) );
  XNOR2_X2 U14488 ( .A(n12426), .B(n12427), .ZN(n12469) );
  OAI21_X4 U14489 ( .B1(n12280), .B2(n12371), .A(n5875), .ZN(n12281) );
  NOR2_X4 U14490 ( .A1(n5044), .A2(n12283), .ZN(n12300) );
  NOR2_X4 U14491 ( .A1(n5044), .A2(n12286), .ZN(n12299) );
  XNOR2_X2 U14492 ( .A(n12302), .B(n4983), .ZN(n12303) );
  NAND2_X2 U14493 ( .A1(aluBoi_multBoi_temppp[59]), .A2(n12304), .ZN(n12305)
         );
  XNOR2_X2 U14494 ( .A(n12306), .B(n12305), .ZN(n12540) );
  INV_X4 U14495 ( .A(n12540), .ZN(n12307) );
  NAND2_X2 U14496 ( .A1(n12528), .A2(n12307), .ZN(net359682) );
  NOR2_X4 U14497 ( .A1(n6438), .A2(n12308), .ZN(aluBoi_multBoi_N67) );
  MUX2_X2 U14498 ( .A(aluBoi_multBoi_temppp[27]), .B(n12309), .S(net367631), 
        .Z(n13679) );
  XOR2_X2 U14499 ( .A(n12311), .B(n12310), .Z(n12313) );
  MUX2_X2 U14500 ( .A(n12313), .B(n12312), .S(net367631), .Z(
        aluBoi_multBoi_N37) );
  XNOR2_X2 U14501 ( .A(n12314), .B(aluBoi_multBoi_temppp[35]), .ZN(n12320) );
  NAND2_X2 U14502 ( .A1(n12316), .A2(n12315), .ZN(n12494) );
  XNOR2_X2 U14503 ( .A(n12317), .B(n5552), .ZN(n12493) );
  NAND2_X2 U14504 ( .A1(n12494), .A2(n12493), .ZN(n12495) );
  NAND2_X2 U14505 ( .A1(n12495), .A2(n12318), .ZN(n12319) );
  XNOR2_X2 U14506 ( .A(n12320), .B(n12319), .ZN(n12321) );
  XNOR2_X2 U14507 ( .A(n12322), .B(net359792), .ZN(n12323) );
  NOR2_X4 U14508 ( .A1(net368481), .A2(n12323), .ZN(aluBoi_multBoi_N45) );
  INV_X4 U14509 ( .A(n12324), .ZN(n12325) );
  INV_X4 U14510 ( .A(net359785), .ZN(net359553) );
  XNOR2_X2 U14511 ( .A(n12328), .B(n12327), .ZN(n12329) );
  XNOR2_X2 U14512 ( .A(n12330), .B(net359540), .ZN(n12331) );
  XNOR2_X2 U14513 ( .A(n12332), .B(n12519), .ZN(n12333) );
  INV_X4 U14514 ( .A(net359767), .ZN(net359512) );
  NAND2_X2 U14515 ( .A1(net359770), .A2(net359771), .ZN(n12334) );
  INV_X4 U14516 ( .A(net359765), .ZN(net359513) );
  INV_X4 U14517 ( .A(net359574), .ZN(net359648) );
  OAI22_X2 U14518 ( .A1(n9729), .A2(net368436), .B1(net368181), .B2(n12342), 
        .ZN(n12447) );
  XNOR2_X2 U14519 ( .A(n12447), .B(n12473), .ZN(n12347) );
  OAI21_X4 U14520 ( .B1(n12345), .B2(n12344), .A(n12568), .ZN(n12461) );
  INV_X4 U14521 ( .A(n12461), .ZN(n12346) );
  OAI21_X4 U14522 ( .B1(n12346), .B2(n12460), .A(n12573), .ZN(n12474) );
  OAI21_X4 U14523 ( .B1(n12352), .B2(n12351), .A(n12350), .ZN(n12356) );
  NAND3_X4 U14524 ( .A1(n12356), .A2(n12427), .A3(n12355), .ZN(n12562) );
  NAND2_X2 U14525 ( .A1(n12357), .A2(n12370), .ZN(n12471) );
  XNOR2_X2 U14526 ( .A(n12426), .B(n12427), .ZN(n12437) );
  NAND2_X2 U14527 ( .A1(n12361), .A2(n5875), .ZN(n12428) );
  INV_X4 U14528 ( .A(n12428), .ZN(n12468) );
  AOI211_X4 U14529 ( .C1(n12362), .C2(n12466), .A(n12468), .B(n12437), .ZN(
        n12366) );
  XNOR2_X2 U14530 ( .A(n12281), .B(n5969), .ZN(n12383) );
  NAND2_X2 U14531 ( .A1(n12378), .A2(n12377), .ZN(n12380) );
  AOI21_X4 U14532 ( .B1(n12389), .B2(n12388), .A(n12387), .ZN(n12390) );
  OAI21_X4 U14533 ( .B1(n5068), .B2(n12397), .A(n12396), .ZN(n12398) );
  NAND4_X2 U14534 ( .A1(net359682), .A2(net359459), .A3(n12538), .A4(net359462), .ZN(n12482) );
  INV_X4 U14535 ( .A(net359681), .ZN(net359680) );
  OAI21_X4 U14536 ( .B1(n12413), .B2(n12414), .A(n12412), .ZN(net359449) );
  OAI221_X2 U14537 ( .B1(net359648), .B2(n12482), .C1(n12417), .C2(n12482), 
        .A(net359650), .ZN(n12488) );
  INV_X4 U14538 ( .A(n12562), .ZN(n12429) );
  INV_X4 U14539 ( .A(n12441), .ZN(n12442) );
  XOR2_X2 U14540 ( .A(n12474), .B(n12473), .Z(n12444) );
  XNOR2_X2 U14541 ( .A(n12445), .B(n12444), .ZN(n12446) );
  NOR2_X4 U14542 ( .A1(n12450), .A2(n12385), .ZN(n12452) );
  OAI21_X4 U14543 ( .B1(n12457), .B2(n12456), .A(n12455), .ZN(n12480) );
  NAND2_X2 U14544 ( .A1(n12461), .A2(n12573), .ZN(n12574) );
  INV_X4 U14545 ( .A(n12473), .ZN(n12570) );
  XNOR2_X2 U14546 ( .A(n12568), .B(n12570), .ZN(n12577) );
  XNOR2_X2 U14547 ( .A(n12574), .B(n12577), .ZN(n12580) );
  NAND2_X2 U14548 ( .A1(n12462), .A2(n12461), .ZN(n12565) );
  OAI21_X4 U14549 ( .B1(n12472), .B2(n12471), .A(n12470), .ZN(n12563) );
  XNOR2_X2 U14550 ( .A(n12474), .B(n12473), .ZN(n12561) );
  NAND2_X2 U14551 ( .A1(n12561), .A2(n12565), .ZN(n12475) );
  XNOR2_X2 U14552 ( .A(n12480), .B(n12559), .ZN(n12543) );
  INV_X4 U14553 ( .A(n6090), .ZN(n12481) );
  OAI221_X2 U14554 ( .B1(n12487), .B2(net377513), .C1(n12487), .C2(net359577), 
        .A(net100619), .ZN(n12486) );
  INV_X4 U14555 ( .A(n12482), .ZN(n12483) );
  OAI211_X2 U14556 ( .C1(n12484), .C2(net359574), .A(n12483), .B(net100619), 
        .ZN(n12485) );
  AOI22_X2 U14557 ( .A1(n12488), .A2(n12487), .B1(n12486), .B2(n12485), .ZN(
        aluBoi_multBoi_N69) );
  XNOR2_X2 U14558 ( .A(n12490), .B(n12489), .ZN(n12492) );
  MUX2_X2 U14559 ( .A(n12492), .B(n12491), .S(net367631), .Z(
        aluBoi_multBoi_N36) );
  INV_X4 U14560 ( .A(n12495), .ZN(n12496) );
  INV_X4 U14561 ( .A(n12500), .ZN(aluBoi_multBoi_N44) );
  INV_X4 U14562 ( .A(n12507), .ZN(aluBoi_multBoi_N56) );
  NAND2_X2 U14563 ( .A1(n12509), .A2(net359537), .ZN(n12513) );
  OAI221_X2 U14564 ( .B1(n12515), .B2(n12514), .C1(n12513), .C2(n12512), .A(
        n12511), .ZN(n12517) );
  NOR2_X4 U14565 ( .A1(net376322), .A2(net359512), .ZN(n12521) );
  NAND3_X4 U14566 ( .A1(n12523), .A2(n12522), .A3(n12521), .ZN(n12525) );
  INV_X4 U14567 ( .A(n12525), .ZN(n12524) );
  XNOR2_X2 U14568 ( .A(n12537), .B(n12536), .ZN(net359475) );
  INV_X4 U14569 ( .A(net359475), .ZN(net359465) );
  INV_X4 U14570 ( .A(net359469), .ZN(net359439) );
  NOR2_X4 U14571 ( .A1(net359451), .A2(n12544), .ZN(n12545) );
  OAI21_X4 U14572 ( .B1(n12546), .B2(n12547), .A(n12545), .ZN(n12556) );
  INV_X4 U14573 ( .A(net359449), .ZN(net359448) );
  XNOR2_X2 U14574 ( .A(n12550), .B(net359418), .ZN(n12553) );
  INV_X4 U14575 ( .A(n12551), .ZN(n12552) );
  AOI21_X4 U14576 ( .B1(n12554), .B2(n12553), .A(n12552), .ZN(n12555) );
  OAI21_X4 U14577 ( .B1(net359439), .B2(n12556), .A(n12555), .ZN(n12591) );
  NAND2_X2 U14578 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  INV_X4 U14579 ( .A(n12567), .ZN(n12581) );
  XNOR2_X2 U14580 ( .A(n12568), .B(n12574), .ZN(n12569) );
  NOR2_X4 U14581 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  NOR2_X4 U14582 ( .A1(n12572), .A2(n12571), .ZN(n12587) );
  INV_X4 U14583 ( .A(n12573), .ZN(n12575) );
  XNOR2_X2 U14584 ( .A(n12576), .B(net359418), .ZN(n12579) );
  XNOR2_X2 U14585 ( .A(n12577), .B(n12583), .ZN(n12578) );
  XNOR2_X2 U14586 ( .A(n12579), .B(n12578), .ZN(n12586) );
  INV_X4 U14587 ( .A(n12580), .ZN(n12582) );
  XNOR2_X2 U14588 ( .A(n12582), .B(n12581), .ZN(n12584) );
  NAND2_X2 U14589 ( .A1(n12584), .A2(n12583), .ZN(n12585) );
  FA_X1 U14590 ( .A(n12587), .B(n12586), .CI(n12585), .S(n12588) );
  XNOR2_X2 U14591 ( .A(n12589), .B(n12588), .ZN(n12590) );
  NAND2_X2 U14592 ( .A1(ifOut_95_), .A2(n6581), .ZN(n12594) );
  NAND2_X2 U14593 ( .A1(idOut_117_), .A2(n6590), .ZN(n12593) );
  NAND2_X2 U14594 ( .A1(n12594), .A2(n12593), .ZN(n4554) );
  NAND2_X2 U14595 ( .A1(n6608), .A2(n5038), .ZN(n13508) );
  XNOR2_X2 U14596 ( .A(iaddr[31]), .B(n9989), .ZN(n12596) );
  NAND2_X2 U14597 ( .A1(n6607), .A2(n5038), .ZN(n13506) );
  NAND2_X2 U14598 ( .A1(ifOut_95_), .A2(n6593), .ZN(n12595) );
  OAI21_X4 U14599 ( .B1(n6601), .B2(n12596), .A(n12595), .ZN(n4555) );
  NAND2_X2 U14600 ( .A1(ifOut_31_), .A2(n6583), .ZN(n12598) );
  NAND2_X2 U14601 ( .A1(n6588), .A2(idOut_70_), .ZN(n12597) );
  NAND2_X2 U14602 ( .A1(n12598), .A2(n12597), .ZN(n4556) );
  NAND2_X2 U14603 ( .A1(n12599), .A2(n12840), .ZN(n12822) );
  INV_X4 U14604 ( .A(n12822), .ZN(n12600) );
  NAND2_X2 U14605 ( .A1(n12800), .A2(iaddr[12]), .ZN(n12799) );
  INV_X4 U14606 ( .A(n12799), .ZN(n12601) );
  NAND2_X2 U14607 ( .A1(n12601), .A2(iaddr[13]), .ZN(n12779) );
  NAND2_X2 U14608 ( .A1(n12781), .A2(iaddr[14]), .ZN(n12780) );
  INV_X4 U14609 ( .A(n12780), .ZN(n12602) );
  NAND2_X2 U14610 ( .A1(n12602), .A2(iaddr[15]), .ZN(n12758) );
  NAND2_X2 U14611 ( .A1(n12760), .A2(iaddr[16]), .ZN(n12759) );
  INV_X4 U14612 ( .A(n12759), .ZN(n12603) );
  NAND2_X2 U14613 ( .A1(n12603), .A2(iaddr[17]), .ZN(n12738) );
  NAND2_X2 U14614 ( .A1(n12740), .A2(iaddr[18]), .ZN(n12739) );
  INV_X4 U14615 ( .A(n12739), .ZN(n12604) );
  NAND2_X2 U14616 ( .A1(n12604), .A2(iaddr[19]), .ZN(n12718) );
  NAND2_X2 U14617 ( .A1(n12720), .A2(iaddr[20]), .ZN(n12719) );
  INV_X4 U14618 ( .A(n12719), .ZN(n12605) );
  NAND2_X2 U14619 ( .A1(n12605), .A2(iaddr[21]), .ZN(n12698) );
  NAND2_X2 U14620 ( .A1(n12700), .A2(iaddr[22]), .ZN(n12699) );
  NAND2_X2 U14621 ( .A1(iaddr[23]), .A2(n12693), .ZN(n12692) );
  NAND2_X2 U14622 ( .A1(n12676), .A2(iaddr[24]), .ZN(n12675) );
  INV_X4 U14623 ( .A(n12675), .ZN(n12606) );
  NAND2_X2 U14624 ( .A1(n12606), .A2(iaddr[25]), .ZN(n12653) );
  NAND2_X2 U14625 ( .A1(n12655), .A2(iaddr[26]), .ZN(n12654) );
  INV_X4 U14626 ( .A(n12654), .ZN(n12607) );
  NAND2_X2 U14627 ( .A1(n12607), .A2(iaddr[27]), .ZN(n12633) );
  NAND2_X2 U14628 ( .A1(n12635), .A2(iaddr[28]), .ZN(n12634) );
  INV_X4 U14629 ( .A(n12634), .ZN(n12608) );
  NAND2_X2 U14630 ( .A1(n12608), .A2(iaddr[29]), .ZN(n12618) );
  NAND2_X2 U14631 ( .A1(iaddr[30]), .A2(n12620), .ZN(n12619) );
  XOR2_X2 U14632 ( .A(n12619), .B(iaddr[31]), .Z(n12610) );
  NAND2_X2 U14633 ( .A1(ifOut_31_), .A2(n6593), .ZN(n12609) );
  NAND2_X2 U14634 ( .A1(ifOut_94_), .A2(n6584), .ZN(n12612) );
  NAND2_X2 U14635 ( .A1(idOut_116_), .A2(n6590), .ZN(n12611) );
  NAND2_X2 U14636 ( .A1(n12612), .A2(n12611), .ZN(n4559) );
  OAI211_X2 U14637 ( .C1(iaddr[30]), .C2(n10010), .A(n12613), .B(n6603), .ZN(
        n12615) );
  NAND2_X2 U14638 ( .A1(ifOut_94_), .A2(n6598), .ZN(n12614) );
  NAND2_X2 U14639 ( .A1(n12615), .A2(n12614), .ZN(n4560) );
  NAND2_X2 U14640 ( .A1(ifOut_30_), .A2(n6584), .ZN(n12617) );
  NAND2_X2 U14641 ( .A1(n6588), .A2(idOut_69_), .ZN(n12616) );
  NAND2_X2 U14642 ( .A1(n12617), .A2(n12616), .ZN(n4561) );
  INV_X4 U14643 ( .A(n12618), .ZN(n12620) );
  OAI211_X2 U14644 ( .C1(iaddr[30]), .C2(n12620), .A(n12619), .B(n6603), .ZN(
        n12622) );
  NAND2_X2 U14645 ( .A1(ifOut_30_), .A2(n6598), .ZN(n12621) );
  NAND2_X2 U14646 ( .A1(n12622), .A2(n12621), .ZN(n4562) );
  NAND2_X2 U14647 ( .A1(ifOut_93_), .A2(n6583), .ZN(n12624) );
  NAND2_X2 U14648 ( .A1(idOut_115_), .A2(n6590), .ZN(n12623) );
  NAND2_X2 U14649 ( .A1(n12624), .A2(n12623), .ZN(n4564) );
  NAND2_X2 U14650 ( .A1(ifOut_93_), .A2(n6598), .ZN(n12626) );
  NAND2_X2 U14651 ( .A1(n12627), .A2(n12626), .ZN(n4565) );
  NAND2_X2 U14652 ( .A1(ifOut_29_), .A2(n6584), .ZN(n12629) );
  NAND2_X2 U14653 ( .A1(n6588), .A2(idOut_68_), .ZN(n12628) );
  NAND2_X2 U14654 ( .A1(n12629), .A2(n12628), .ZN(n4566) );
  XNOR2_X2 U14655 ( .A(n12634), .B(n5571), .ZN(n12630) );
  OAI22_X2 U14656 ( .A1(n6601), .A2(n12630), .B1(n6594), .B2(n5599), .ZN(n4567) );
  NAND2_X2 U14657 ( .A1(ifOut_28_), .A2(n6584), .ZN(n12632) );
  NAND2_X2 U14658 ( .A1(n6588), .A2(idOut_67_), .ZN(n12631) );
  NAND2_X2 U14659 ( .A1(n12632), .A2(n12631), .ZN(n4569) );
  INV_X4 U14660 ( .A(n12633), .ZN(n12635) );
  OAI211_X2 U14661 ( .C1(iaddr[28]), .C2(n12635), .A(n12634), .B(n6603), .ZN(
        n12637) );
  NAND2_X2 U14662 ( .A1(ifOut_28_), .A2(n6598), .ZN(n12636) );
  NAND2_X2 U14663 ( .A1(n12637), .A2(n12636), .ZN(n4570) );
  NAND2_X2 U14664 ( .A1(ifOut_92_), .A2(n6584), .ZN(n12639) );
  NAND2_X2 U14665 ( .A1(idOut_114_), .A2(n6590), .ZN(n12638) );
  NAND2_X2 U14666 ( .A1(n12639), .A2(n12638), .ZN(n4571) );
  NAND2_X2 U14667 ( .A1(ifOut_92_), .A2(n6598), .ZN(n12641) );
  NAND2_X2 U14668 ( .A1(n12642), .A2(n12641), .ZN(n4572) );
  NAND2_X2 U14669 ( .A1(ifOut_91_), .A2(n6584), .ZN(n12644) );
  NAND2_X2 U14670 ( .A1(idOut_113_), .A2(n6589), .ZN(n12643) );
  NAND2_X2 U14671 ( .A1(n12644), .A2(n12643), .ZN(n4574) );
  NAND2_X2 U14672 ( .A1(ifOut_91_), .A2(n6598), .ZN(n12646) );
  NAND2_X2 U14673 ( .A1(n12647), .A2(n12646), .ZN(n4575) );
  NAND2_X2 U14674 ( .A1(ifOut_27_), .A2(n6584), .ZN(n12649) );
  NAND2_X2 U14675 ( .A1(n6588), .A2(idOut_66_), .ZN(n12648) );
  NAND2_X2 U14676 ( .A1(n12649), .A2(n12648), .ZN(n4576) );
  XNOR2_X2 U14677 ( .A(n12654), .B(n5580), .ZN(n12650) );
  OAI22_X2 U14678 ( .A1(n6601), .A2(n12650), .B1(n6597), .B2(n5600), .ZN(n4577) );
  NAND2_X2 U14679 ( .A1(ifOut_26_), .A2(n6584), .ZN(n12652) );
  NAND2_X2 U14680 ( .A1(n6588), .A2(idOut_65_), .ZN(n12651) );
  NAND2_X2 U14681 ( .A1(n12652), .A2(n12651), .ZN(n4579) );
  INV_X4 U14682 ( .A(n12653), .ZN(n12655) );
  OAI211_X2 U14683 ( .C1(iaddr[26]), .C2(n12655), .A(n12654), .B(n6603), .ZN(
        n12657) );
  NAND2_X2 U14684 ( .A1(ifOut_26_), .A2(n6598), .ZN(n12656) );
  NAND2_X2 U14685 ( .A1(n12657), .A2(n12656), .ZN(n4580) );
  NAND2_X2 U14686 ( .A1(ifOut_90_), .A2(n6584), .ZN(n12659) );
  NAND2_X2 U14687 ( .A1(idOut_112_), .A2(n6589), .ZN(n12658) );
  NAND2_X2 U14688 ( .A1(n12659), .A2(n12658), .ZN(n4581) );
  INV_X4 U14689 ( .A(n12666), .ZN(n12661) );
  OAI211_X2 U14690 ( .C1(iaddr[26]), .C2(n12661), .A(n12660), .B(n6603), .ZN(
        n12663) );
  NAND2_X2 U14691 ( .A1(ifOut_90_), .A2(n6598), .ZN(n12662) );
  NAND2_X2 U14692 ( .A1(n12663), .A2(n12662), .ZN(n4582) );
  NAND2_X2 U14693 ( .A1(ifOut_89_), .A2(n6584), .ZN(n12665) );
  NAND2_X2 U14694 ( .A1(idOut_111_), .A2(n6590), .ZN(n12664) );
  NAND2_X2 U14695 ( .A1(n12665), .A2(n12664), .ZN(n4584) );
  OAI211_X2 U14696 ( .C1(iaddr[25]), .C2(n12667), .A(n12666), .B(n6603), .ZN(
        n12669) );
  NAND2_X2 U14697 ( .A1(ifOut_89_), .A2(n6598), .ZN(n12668) );
  NAND2_X2 U14698 ( .A1(n12669), .A2(n12668), .ZN(n4585) );
  NAND2_X2 U14699 ( .A1(ifOut_25_), .A2(n6584), .ZN(n12671) );
  NAND2_X2 U14700 ( .A1(n6590), .A2(idOut_64_), .ZN(n12670) );
  NAND2_X2 U14701 ( .A1(n12671), .A2(n12670), .ZN(n4586) );
  XOR2_X2 U14702 ( .A(n12675), .B(iaddr[25]), .Z(n12672) );
  OAI22_X2 U14703 ( .A1(n6601), .A2(n12672), .B1(n6597), .B2(n5601), .ZN(n4587) );
  NAND2_X2 U14704 ( .A1(ifOut_24_), .A2(n6584), .ZN(n12674) );
  NAND2_X2 U14705 ( .A1(n6588), .A2(idOut_63_), .ZN(n12673) );
  NAND2_X2 U14706 ( .A1(n12674), .A2(n12673), .ZN(n4589) );
  INV_X4 U14707 ( .A(n12692), .ZN(n12676) );
  OAI211_X2 U14708 ( .C1(iaddr[24]), .C2(n12676), .A(n12675), .B(n6603), .ZN(
        n12678) );
  NAND2_X2 U14709 ( .A1(ifOut_24_), .A2(n6598), .ZN(n12677) );
  NAND2_X2 U14710 ( .A1(n12678), .A2(n12677), .ZN(n4590) );
  NAND2_X2 U14711 ( .A1(ifOut_88_), .A2(n6584), .ZN(n12680) );
  NAND2_X2 U14712 ( .A1(idOut_110_), .A2(n6589), .ZN(n12679) );
  NAND2_X2 U14713 ( .A1(n12680), .A2(n12679), .ZN(n4591) );
  OAI211_X2 U14714 ( .C1(iaddr[24]), .C2(n12682), .A(n12681), .B(n6603), .ZN(
        n12684) );
  NAND2_X2 U14715 ( .A1(ifOut_88_), .A2(n6598), .ZN(n12683) );
  NAND2_X2 U14716 ( .A1(n12684), .A2(n12683), .ZN(n4592) );
  NAND2_X2 U14717 ( .A1(ifOut_87_), .A2(n6584), .ZN(n12686) );
  NAND2_X2 U14718 ( .A1(idOut_109_), .A2(n6589), .ZN(n12685) );
  NAND2_X2 U14719 ( .A1(n12686), .A2(n12685), .ZN(n4594) );
  NAND2_X2 U14720 ( .A1(ifOut_87_), .A2(n6598), .ZN(n12688) );
  NAND2_X2 U14721 ( .A1(n12689), .A2(n12688), .ZN(n4595) );
  NAND2_X2 U14722 ( .A1(ifOut_23_), .A2(n6584), .ZN(n12691) );
  NAND2_X2 U14723 ( .A1(n6588), .A2(idOut_62_), .ZN(n12690) );
  NAND2_X2 U14724 ( .A1(n12691), .A2(n12690), .ZN(n4596) );
  INV_X4 U14725 ( .A(n12699), .ZN(n12693) );
  OAI211_X2 U14726 ( .C1(iaddr[23]), .C2(n12693), .A(n12692), .B(n6603), .ZN(
        n12695) );
  NAND2_X2 U14727 ( .A1(ifOut_23_), .A2(n6598), .ZN(n12694) );
  NAND2_X2 U14728 ( .A1(n12695), .A2(n12694), .ZN(n4597) );
  NAND2_X2 U14729 ( .A1(ifOut_22_), .A2(n6584), .ZN(n12697) );
  NAND2_X2 U14730 ( .A1(n6588), .A2(idOut_61_), .ZN(n12696) );
  NAND2_X2 U14731 ( .A1(n12697), .A2(n12696), .ZN(n4599) );
  INV_X4 U14732 ( .A(n12698), .ZN(n12700) );
  OAI211_X2 U14733 ( .C1(iaddr[22]), .C2(n12700), .A(n12699), .B(n6603), .ZN(
        n12702) );
  NAND2_X2 U14734 ( .A1(ifOut_22_), .A2(n6598), .ZN(n12701) );
  NAND2_X2 U14735 ( .A1(n12702), .A2(n12701), .ZN(n4600) );
  NAND2_X2 U14736 ( .A1(ifOut_86_), .A2(n6584), .ZN(n12704) );
  NAND2_X2 U14737 ( .A1(idOut_108_), .A2(n6589), .ZN(n12703) );
  NAND2_X2 U14738 ( .A1(n12704), .A2(n12703), .ZN(n4601) );
  NAND2_X2 U14739 ( .A1(ifOut_86_), .A2(n6598), .ZN(n12706) );
  NAND2_X2 U14740 ( .A1(n12707), .A2(n12706), .ZN(n4602) );
  NAND2_X2 U14741 ( .A1(ifOut_85_), .A2(n6584), .ZN(n12709) );
  NAND2_X2 U14742 ( .A1(idOut_107_), .A2(n6589), .ZN(n12708) );
  NAND2_X2 U14743 ( .A1(n12709), .A2(n12708), .ZN(n4604) );
  OAI211_X2 U14744 ( .C1(iaddr[21]), .C2(n10144), .A(n12710), .B(n6603), .ZN(
        n12712) );
  NAND2_X2 U14745 ( .A1(ifOut_85_), .A2(n6598), .ZN(n12711) );
  NAND2_X2 U14746 ( .A1(n12712), .A2(n12711), .ZN(n4605) );
  NAND2_X2 U14747 ( .A1(ifOut_21_), .A2(n6584), .ZN(n12714) );
  NAND2_X2 U14748 ( .A1(n6590), .A2(idOut_60_), .ZN(n12713) );
  NAND2_X2 U14749 ( .A1(n12714), .A2(n12713), .ZN(n4606) );
  XNOR2_X2 U14750 ( .A(n12719), .B(n5562), .ZN(n12715) );
  OAI22_X2 U14751 ( .A1(n6601), .A2(n12715), .B1(n6597), .B2(n5602), .ZN(n4607) );
  NAND2_X2 U14752 ( .A1(ifOut_20_), .A2(n6584), .ZN(n12717) );
  NAND2_X2 U14753 ( .A1(n6588), .A2(idOut_59_), .ZN(n12716) );
  NAND2_X2 U14754 ( .A1(n12717), .A2(n12716), .ZN(n4609) );
  INV_X4 U14755 ( .A(n12718), .ZN(n12720) );
  OAI211_X2 U14756 ( .C1(iaddr[20]), .C2(n12720), .A(n12719), .B(n6603), .ZN(
        n12722) );
  NAND2_X2 U14757 ( .A1(ifOut_20_), .A2(n6598), .ZN(n12721) );
  NAND2_X2 U14758 ( .A1(n12722), .A2(n12721), .ZN(n4610) );
  NAND2_X2 U14759 ( .A1(ifOut_84_), .A2(n6584), .ZN(n12724) );
  NAND2_X2 U14760 ( .A1(idOut_106_), .A2(n6589), .ZN(n12723) );
  NAND2_X2 U14761 ( .A1(n12724), .A2(n12723), .ZN(n4611) );
  OAI211_X2 U14762 ( .C1(iaddr[20]), .C2(n10156), .A(n12725), .B(n6603), .ZN(
        n12727) );
  NAND2_X2 U14763 ( .A1(ifOut_84_), .A2(n6598), .ZN(n12726) );
  NAND2_X2 U14764 ( .A1(n12727), .A2(n12726), .ZN(n4612) );
  NAND2_X2 U14765 ( .A1(ifOut_83_), .A2(n6584), .ZN(n12729) );
  NAND2_X2 U14766 ( .A1(idOut_105_), .A2(n6589), .ZN(n12728) );
  NAND2_X2 U14767 ( .A1(n12729), .A2(n12728), .ZN(n4614) );
  OAI211_X2 U14768 ( .C1(iaddr[19]), .C2(n10161), .A(n12730), .B(n6603), .ZN(
        n12732) );
  NAND2_X2 U14769 ( .A1(ifOut_83_), .A2(n6598), .ZN(n12731) );
  NAND2_X2 U14770 ( .A1(n12732), .A2(n12731), .ZN(n4615) );
  NAND2_X2 U14771 ( .A1(ifOut_19_), .A2(n6584), .ZN(n12734) );
  NAND2_X2 U14772 ( .A1(n6588), .A2(idOut_58_), .ZN(n12733) );
  NAND2_X2 U14773 ( .A1(n12734), .A2(n12733), .ZN(n4616) );
  XNOR2_X2 U14774 ( .A(n12739), .B(n5563), .ZN(n12735) );
  OAI22_X2 U14775 ( .A1(n6601), .A2(n12735), .B1(n6597), .B2(n5603), .ZN(n4617) );
  NAND2_X2 U14776 ( .A1(ifOut_18_), .A2(n6584), .ZN(n12737) );
  NAND2_X2 U14777 ( .A1(n6588), .A2(idOut_57_), .ZN(n12736) );
  NAND2_X2 U14778 ( .A1(n12737), .A2(n12736), .ZN(n4619) );
  INV_X4 U14779 ( .A(n12738), .ZN(n12740) );
  OAI211_X2 U14780 ( .C1(iaddr[18]), .C2(n12740), .A(n12739), .B(n6603), .ZN(
        n12742) );
  NAND2_X2 U14781 ( .A1(ifOut_18_), .A2(n6598), .ZN(n12741) );
  NAND2_X2 U14782 ( .A1(n12742), .A2(n12741), .ZN(n4620) );
  NAND2_X2 U14783 ( .A1(ifOut_82_), .A2(n6584), .ZN(n12744) );
  NAND2_X2 U14784 ( .A1(idOut_104_), .A2(n6589), .ZN(n12743) );
  NAND2_X2 U14785 ( .A1(n12744), .A2(n12743), .ZN(n4621) );
  OAI211_X2 U14786 ( .C1(iaddr[18]), .C2(n10181), .A(n12745), .B(n6603), .ZN(
        n12747) );
  NAND2_X2 U14787 ( .A1(ifOut_82_), .A2(n6598), .ZN(n12746) );
  NAND2_X2 U14788 ( .A1(n12747), .A2(n12746), .ZN(n4622) );
  NAND2_X2 U14789 ( .A1(ifOut_81_), .A2(n6584), .ZN(n12749) );
  NAND2_X2 U14790 ( .A1(idOut_103_), .A2(n6589), .ZN(n12748) );
  NAND2_X2 U14791 ( .A1(n12749), .A2(n12748), .ZN(n4624) );
  NAND2_X2 U14792 ( .A1(ifOut_81_), .A2(n6598), .ZN(n12751) );
  NAND2_X2 U14793 ( .A1(n12752), .A2(n12751), .ZN(n4625) );
  NAND2_X2 U14794 ( .A1(ifOut_17_), .A2(n6584), .ZN(n12754) );
  NAND2_X2 U14795 ( .A1(n6588), .A2(idOut_56_), .ZN(n12753) );
  NAND2_X2 U14796 ( .A1(n12754), .A2(n12753), .ZN(n4626) );
  XNOR2_X2 U14797 ( .A(n12759), .B(n5581), .ZN(n12755) );
  OAI22_X2 U14798 ( .A1(n6601), .A2(n12755), .B1(n6597), .B2(n5604), .ZN(n4627) );
  NAND2_X2 U14799 ( .A1(ifOut_16_), .A2(n6583), .ZN(n12757) );
  NAND2_X2 U14800 ( .A1(n6588), .A2(idOut_55_), .ZN(n12756) );
  NAND2_X2 U14801 ( .A1(n12757), .A2(n12756), .ZN(n4629) );
  INV_X4 U14802 ( .A(n12758), .ZN(n12760) );
  OAI211_X2 U14803 ( .C1(iaddr[16]), .C2(n12760), .A(n12759), .B(n6603), .ZN(
        n12762) );
  NAND2_X2 U14804 ( .A1(ifOut_16_), .A2(n6598), .ZN(n12761) );
  NAND2_X2 U14805 ( .A1(n12762), .A2(n12761), .ZN(n4630) );
  NAND2_X2 U14806 ( .A1(ifOut_80_), .A2(n6583), .ZN(n12764) );
  NAND2_X2 U14807 ( .A1(idOut_102_), .A2(n6589), .ZN(n12763) );
  NAND2_X2 U14808 ( .A1(n12764), .A2(n12763), .ZN(n4631) );
  NAND2_X2 U14809 ( .A1(ifOut_80_), .A2(n6598), .ZN(n12766) );
  NAND2_X2 U14810 ( .A1(n12767), .A2(n12766), .ZN(n4632) );
  NAND2_X2 U14811 ( .A1(ifOut_79_), .A2(n6583), .ZN(n12769) );
  NAND2_X2 U14812 ( .A1(idOut_101_), .A2(n6588), .ZN(n12768) );
  NAND2_X2 U14813 ( .A1(n12769), .A2(n12768), .ZN(n13609) );
  OAI211_X2 U14814 ( .C1(iaddr[15]), .C2(n12771), .A(n12770), .B(n6603), .ZN(
        n12773) );
  NAND2_X2 U14815 ( .A1(ifOut_79_), .A2(n6598), .ZN(n12772) );
  NAND2_X2 U14816 ( .A1(n12773), .A2(n12772), .ZN(n4635) );
  NAND2_X2 U14817 ( .A1(ifOut_15_), .A2(n6583), .ZN(n12775) );
  NAND2_X2 U14818 ( .A1(idOut_54_), .A2(n6589), .ZN(n12774) );
  NAND2_X2 U14819 ( .A1(n12775), .A2(n12774), .ZN(n4636) );
  XNOR2_X2 U14820 ( .A(n12780), .B(n5574), .ZN(n12776) );
  OAI22_X2 U14821 ( .A1(n6601), .A2(n12776), .B1(n6596), .B2(n5605), .ZN(n4637) );
  NAND2_X2 U14822 ( .A1(ifOut_14_), .A2(n6583), .ZN(n12778) );
  NAND2_X2 U14823 ( .A1(idOut_53_), .A2(n6588), .ZN(n12777) );
  NAND2_X2 U14824 ( .A1(n12778), .A2(n12777), .ZN(n4639) );
  INV_X4 U14825 ( .A(n12779), .ZN(n12781) );
  OAI211_X2 U14826 ( .C1(iaddr[14]), .C2(n12781), .A(n12780), .B(n6603), .ZN(
        n12783) );
  NAND2_X2 U14827 ( .A1(ifOut_14_), .A2(n6598), .ZN(n12782) );
  NAND2_X2 U14828 ( .A1(n12783), .A2(n12782), .ZN(n4640) );
  NAND2_X2 U14829 ( .A1(ifOut_78_), .A2(n6583), .ZN(n12785) );
  NAND2_X2 U14830 ( .A1(idOut_100_), .A2(n6588), .ZN(n12784) );
  NAND2_X2 U14831 ( .A1(n12785), .A2(n12784), .ZN(n4641) );
  OAI211_X2 U14832 ( .C1(iaddr[14]), .C2(n10234), .A(n12786), .B(n6603), .ZN(
        n12788) );
  NAND2_X2 U14833 ( .A1(ifOut_78_), .A2(n6598), .ZN(n12787) );
  NAND2_X2 U14834 ( .A1(n12788), .A2(n12787), .ZN(n4642) );
  NAND2_X2 U14835 ( .A1(ifOut_77_), .A2(n6583), .ZN(n12790) );
  NAND2_X2 U14836 ( .A1(idOut_99_), .A2(n6589), .ZN(n12789) );
  NAND2_X2 U14837 ( .A1(n12790), .A2(n12789), .ZN(n13628) );
  OAI211_X2 U14838 ( .C1(iaddr[13]), .C2(n10239), .A(n12791), .B(n6603), .ZN(
        n12793) );
  NAND2_X2 U14839 ( .A1(ifOut_77_), .A2(n6598), .ZN(n12792) );
  NAND2_X2 U14840 ( .A1(n12793), .A2(n12792), .ZN(n4645) );
  NAND2_X2 U14841 ( .A1(ifOut_13_), .A2(n6583), .ZN(n12795) );
  NAND2_X2 U14842 ( .A1(idOut_52_), .A2(n6588), .ZN(n12794) );
  NAND2_X2 U14843 ( .A1(n12795), .A2(n12794), .ZN(n4646) );
  XNOR2_X2 U14844 ( .A(n12799), .B(n5564), .ZN(n12796) );
  OAI22_X2 U14845 ( .A1(n6601), .A2(n12796), .B1(n6596), .B2(n5606), .ZN(n4647) );
  NAND2_X2 U14846 ( .A1(ifOut_12_), .A2(n6583), .ZN(n12798) );
  NAND2_X2 U14847 ( .A1(idOut_51_), .A2(n6588), .ZN(n12797) );
  NAND2_X2 U14848 ( .A1(n12798), .A2(n12797), .ZN(n4649) );
  INV_X4 U14849 ( .A(n12816), .ZN(n12800) );
  OAI211_X2 U14850 ( .C1(iaddr[12]), .C2(n12800), .A(n12799), .B(n6603), .ZN(
        n12802) );
  NAND2_X2 U14851 ( .A1(ifOut_12_), .A2(n6598), .ZN(n12801) );
  NAND2_X2 U14852 ( .A1(n12802), .A2(n12801), .ZN(n4650) );
  NAND2_X2 U14853 ( .A1(ifOut_76_), .A2(n6583), .ZN(n12804) );
  NAND2_X2 U14854 ( .A1(idOut_98_), .A2(n6589), .ZN(n12803) );
  NAND2_X2 U14855 ( .A1(n12804), .A2(n12803), .ZN(n4651) );
  OAI211_X2 U14856 ( .C1(iaddr[12]), .C2(n10259), .A(n12805), .B(n6603), .ZN(
        n12807) );
  NAND2_X2 U14857 ( .A1(ifOut_76_), .A2(n6598), .ZN(n12806) );
  NAND2_X2 U14858 ( .A1(n12807), .A2(n12806), .ZN(n4652) );
  NAND2_X2 U14859 ( .A1(ifOut_75_), .A2(n6583), .ZN(n12809) );
  NAND2_X2 U14860 ( .A1(idOut_97_), .A2(n6588), .ZN(n12808) );
  NAND2_X2 U14861 ( .A1(n12809), .A2(n12808), .ZN(n13627) );
  NAND2_X2 U14862 ( .A1(ifOut_75_), .A2(n6598), .ZN(n12812) );
  NAND2_X2 U14863 ( .A1(n12813), .A2(n12812), .ZN(n4655) );
  NAND2_X2 U14864 ( .A1(ifOut_11_), .A2(n6583), .ZN(n12815) );
  NAND2_X2 U14865 ( .A1(idOut_50_), .A2(n6588), .ZN(n12814) );
  NAND2_X2 U14866 ( .A1(n12815), .A2(n12814), .ZN(n4656) );
  OAI211_X2 U14867 ( .C1(n12817), .C2(iaddr[11]), .A(n12816), .B(n6603), .ZN(
        n12819) );
  NAND2_X2 U14868 ( .A1(ifOut_11_), .A2(n6598), .ZN(n12818) );
  NAND2_X2 U14869 ( .A1(n12819), .A2(n12818), .ZN(n4657) );
  NAND2_X2 U14870 ( .A1(ifOut_10_), .A2(n6583), .ZN(n12821) );
  NAND2_X2 U14871 ( .A1(idOut_49_), .A2(n6589), .ZN(n12820) );
  NAND2_X2 U14872 ( .A1(n12821), .A2(n12820), .ZN(n13611) );
  XNOR2_X2 U14873 ( .A(n12822), .B(n5478), .ZN(n12823) );
  OAI22_X2 U14874 ( .A1(n6601), .A2(n12823), .B1(n6596), .B2(n5607), .ZN(n4660) );
  NAND2_X2 U14875 ( .A1(ifOut_74_), .A2(n6583), .ZN(n12825) );
  NAND2_X2 U14876 ( .A1(idOut_96_), .A2(n6588), .ZN(n12824) );
  NAND2_X2 U14877 ( .A1(n12825), .A2(n12824), .ZN(n4661) );
  XNOR2_X2 U14878 ( .A(n12826), .B(n5478), .ZN(n12827) );
  OAI22_X2 U14879 ( .A1(n6601), .A2(n12827), .B1(n6596), .B2(n5489), .ZN(n4662) );
  NAND2_X2 U14880 ( .A1(ifOut_73_), .A2(n6583), .ZN(n12829) );
  NAND2_X2 U14881 ( .A1(idOut_95_), .A2(n6588), .ZN(n12828) );
  NAND2_X2 U14882 ( .A1(n12829), .A2(n12828), .ZN(n13626) );
  NAND2_X2 U14883 ( .A1(iaddr[9]), .A2(n6603), .ZN(n12842) );
  INV_X4 U14884 ( .A(n12842), .ZN(n12831) );
  NAND2_X2 U14885 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  INV_X4 U14886 ( .A(n12832), .ZN(n12839) );
  INV_X4 U14887 ( .A(n12833), .ZN(n12834) );
  NAND2_X2 U14888 ( .A1(n12834), .A2(n6603), .ZN(n12841) );
  MUX2_X2 U14889 ( .A(n12842), .B(n12841), .S(n5347), .Z(n12835) );
  NAND2_X2 U14890 ( .A1(n12836), .A2(n12835), .ZN(n4665) );
  NAND2_X2 U14891 ( .A1(ifOut_9_), .A2(n6583), .ZN(n12838) );
  NAND2_X2 U14892 ( .A1(idOut_48_), .A2(n6588), .ZN(n12837) );
  NAND2_X2 U14893 ( .A1(n12838), .A2(n12837), .ZN(n13610) );
  MUX2_X2 U14894 ( .A(n12842), .B(n12841), .S(n12840), .Z(n12843) );
  NAND2_X2 U14895 ( .A1(n12844), .A2(n12843), .ZN(n4667) );
  NAND2_X2 U14896 ( .A1(ifOut_72_), .A2(n6583), .ZN(n12846) );
  NAND2_X2 U14897 ( .A1(idOut_94_), .A2(n6588), .ZN(n12845) );
  NAND2_X2 U14898 ( .A1(n12846), .A2(n12845), .ZN(n4669) );
  XOR2_X2 U14899 ( .A(n12854), .B(iaddr[8]), .Z(n12847) );
  OAI22_X2 U14900 ( .A1(n6601), .A2(n12847), .B1(n6596), .B2(n5506), .ZN(n4670) );
  NAND2_X2 U14901 ( .A1(ifOut_8_), .A2(n6583), .ZN(n12849) );
  NAND2_X2 U14902 ( .A1(idOut_47_), .A2(n6588), .ZN(n12848) );
  NAND2_X2 U14903 ( .A1(n12849), .A2(n12848), .ZN(n4671) );
  XOR2_X2 U14904 ( .A(iaddr[8]), .B(n12859), .Z(n12850) );
  OAI22_X2 U14905 ( .A1(n6601), .A2(n12850), .B1(n6596), .B2(n5608), .ZN(n4672) );
  NAND2_X2 U14906 ( .A1(ifOut_71_), .A2(n6583), .ZN(n12852) );
  NAND2_X2 U14907 ( .A1(idOut_93_), .A2(n6588), .ZN(n12851) );
  NAND2_X2 U14908 ( .A1(n12852), .A2(n12851), .ZN(n13625) );
  NAND2_X2 U14909 ( .A1(ifOut_71_), .A2(n6598), .ZN(n12855) );
  NAND2_X2 U14910 ( .A1(n12856), .A2(n12855), .ZN(n4675) );
  NAND2_X2 U14911 ( .A1(ifOut_7_), .A2(n6583), .ZN(n12858) );
  NAND2_X2 U14912 ( .A1(idOut_46_), .A2(n6588), .ZN(n12857) );
  NAND2_X2 U14913 ( .A1(n12858), .A2(n12857), .ZN(n4676) );
  NAND2_X2 U14914 ( .A1(ifOut_7_), .A2(n6598), .ZN(n12860) );
  NAND2_X2 U14915 ( .A1(n12861), .A2(n12860), .ZN(n4677) );
  NAND2_X2 U14916 ( .A1(ifOut_70_), .A2(n6583), .ZN(n12863) );
  NAND2_X2 U14917 ( .A1(idOut_92_), .A2(n6590), .ZN(n12862) );
  NAND2_X2 U14918 ( .A1(n12863), .A2(n12862), .ZN(n4679) );
  XOR2_X2 U14919 ( .A(n12870), .B(iaddr[6]), .Z(n12864) );
  OAI22_X2 U14920 ( .A1(n6601), .A2(n12864), .B1(n6596), .B2(n5490), .ZN(n4680) );
  NAND2_X2 U14921 ( .A1(ifOut_6_), .A2(n6583), .ZN(n12866) );
  NAND2_X2 U14922 ( .A1(n6590), .A2(idOut_45_), .ZN(n12865) );
  NAND2_X2 U14923 ( .A1(n12866), .A2(n12865), .ZN(n4681) );
  XNOR2_X2 U14924 ( .A(iaddr[6]), .B(n12875), .ZN(n12867) );
  OAI22_X2 U14925 ( .A1(n6601), .A2(n12867), .B1(n6596), .B2(n5609), .ZN(n4682) );
  NAND2_X2 U14926 ( .A1(ifOut_69_), .A2(n6583), .ZN(n12869) );
  NAND2_X2 U14927 ( .A1(idOut_91_), .A2(n6588), .ZN(n12868) );
  NAND2_X2 U14928 ( .A1(n12869), .A2(n12868), .ZN(n13624) );
  OAI211_X2 U14929 ( .C1(iaddr[5]), .C2(n5347), .A(n12870), .B(n6604), .ZN(
        n12872) );
  NAND2_X2 U14930 ( .A1(ifOut_69_), .A2(n6598), .ZN(n12871) );
  NAND2_X2 U14931 ( .A1(n12872), .A2(n12871), .ZN(n4685) );
  NAND2_X2 U14932 ( .A1(ifOut_5_), .A2(n6583), .ZN(n12874) );
  NAND2_X2 U14933 ( .A1(n6588), .A2(idOut_44_), .ZN(n12873) );
  NAND2_X2 U14934 ( .A1(n12874), .A2(n12873), .ZN(n4686) );
  INV_X4 U14935 ( .A(n12875), .ZN(n12878) );
  NAND2_X2 U14936 ( .A1(n12876), .A2(n5509), .ZN(n12877) );
  NAND2_X2 U14937 ( .A1(ifOut_5_), .A2(n6598), .ZN(n12879) );
  NAND2_X2 U14938 ( .A1(n12880), .A2(n12879), .ZN(n4687) );
  NAND2_X2 U14939 ( .A1(ifOut_68_), .A2(n6582), .ZN(n12882) );
  NAND2_X2 U14940 ( .A1(idOut_90_), .A2(n6588), .ZN(n12881) );
  NAND2_X2 U14941 ( .A1(n12882), .A2(n12881), .ZN(n4689) );
  XOR2_X2 U14942 ( .A(n12883), .B(iaddr[4]), .Z(n12884) );
  OAI22_X2 U14943 ( .A1(n6601), .A2(n12884), .B1(n6596), .B2(n5507), .ZN(n4690) );
  NAND2_X2 U14944 ( .A1(ifOut_4_), .A2(n6582), .ZN(n12886) );
  NAND2_X2 U14945 ( .A1(n6588), .A2(idOut_43_), .ZN(n12885) );
  NAND2_X2 U14946 ( .A1(n12886), .A2(n12885), .ZN(n4691) );
  NAND2_X2 U14947 ( .A1(ifOut_4_), .A2(n6598), .ZN(n12888) );
  NAND2_X2 U14948 ( .A1(n6603), .A2(n5477), .ZN(n12897) );
  MUX2_X2 U14949 ( .A(n12891), .B(n12897), .S(iaddr[4]), .Z(n12887) );
  NAND2_X2 U14950 ( .A1(n12888), .A2(n12887), .ZN(n4692) );
  NAND2_X2 U14951 ( .A1(ifOut_67_), .A2(n6582), .ZN(n12890) );
  NAND2_X2 U14952 ( .A1(idOut_89_), .A2(n6588), .ZN(n12889) );
  NAND2_X2 U14953 ( .A1(n12890), .A2(n12889), .ZN(n13623) );
  NAND2_X2 U14954 ( .A1(ifOut_67_), .A2(n6598), .ZN(n12893) );
  MUX2_X2 U14955 ( .A(n12891), .B(n12897), .S(iaddr[2]), .Z(n12892) );
  NAND2_X2 U14956 ( .A1(n12893), .A2(n12892), .ZN(n4695) );
  NAND2_X2 U14957 ( .A1(ifOut_3_), .A2(n6582), .ZN(n12895) );
  NAND2_X2 U14958 ( .A1(n6587), .A2(idOut_42_), .ZN(n12894) );
  NAND2_X2 U14959 ( .A1(n12895), .A2(n12894), .ZN(n4696) );
  NAND2_X2 U14960 ( .A1(ifOut_3_), .A2(n6598), .ZN(n12896) );
  NAND2_X2 U14961 ( .A1(n12897), .A2(n12896), .ZN(n4697) );
  NAND2_X2 U14962 ( .A1(ifOut_2_), .A2(n6582), .ZN(n12899) );
  NAND2_X2 U14963 ( .A1(n6587), .A2(idOut_41_), .ZN(n12898) );
  NAND2_X2 U14964 ( .A1(n12899), .A2(n12898), .ZN(n4699) );
  OAI22_X2 U14965 ( .A1(n6601), .A2(n5355), .B1(n6596), .B2(n5610), .ZN(n4700)
         );
  NAND2_X2 U14966 ( .A1(ifOut_66_), .A2(n6582), .ZN(n12901) );
  NAND2_X2 U14967 ( .A1(n12901), .A2(n12900), .ZN(n4701) );
  OAI22_X2 U14968 ( .A1(iaddr[2]), .A2(n6602), .B1(n6596), .B2(n5508), .ZN(
        n4702) );
  NAND2_X2 U14969 ( .A1(ifOut_1_), .A2(n6582), .ZN(n12903) );
  NAND2_X2 U14970 ( .A1(n6587), .A2(idOut_40_), .ZN(n12902) );
  NAND2_X2 U14971 ( .A1(n12903), .A2(n12902), .ZN(n4704) );
  NAND2_X2 U14972 ( .A1(iaddr[1]), .A2(n6604), .ZN(n12908) );
  NAND2_X2 U14973 ( .A1(ifOut_1_), .A2(n6593), .ZN(n12904) );
  NAND2_X2 U14974 ( .A1(n12908), .A2(n12904), .ZN(n4705) );
  NAND2_X2 U14975 ( .A1(idOut_87_), .A2(n6588), .ZN(n12905) );
  NAND2_X2 U14976 ( .A1(n12906), .A2(n12905), .ZN(n4706) );
  NAND2_X2 U14977 ( .A1(ifOut_65_), .A2(n6593), .ZN(n12907) );
  NAND2_X2 U14978 ( .A1(n12908), .A2(n12907), .ZN(n4707) );
  NAND2_X2 U14979 ( .A1(ifOut_0_), .A2(n6582), .ZN(n12910) );
  NAND2_X2 U14980 ( .A1(n6587), .A2(idOut_39_), .ZN(n12909) );
  NAND2_X2 U14981 ( .A1(n12910), .A2(n12909), .ZN(n4709) );
  NAND2_X2 U14982 ( .A1(iaddr[0]), .A2(n6604), .ZN(n12915) );
  NAND2_X2 U14983 ( .A1(ifOut_0_), .A2(n6593), .ZN(n12911) );
  NAND2_X2 U14984 ( .A1(n12915), .A2(n12911), .ZN(n4710) );
  NAND2_X2 U14985 ( .A1(ifOut_64_), .A2(n6582), .ZN(n12913) );
  NAND2_X2 U14986 ( .A1(idOut_86_), .A2(n6588), .ZN(n12912) );
  NAND2_X2 U14987 ( .A1(n12913), .A2(n12912), .ZN(n4711) );
  NAND2_X2 U14988 ( .A1(ifOut_64_), .A2(n6598), .ZN(n12914) );
  NAND2_X2 U14989 ( .A1(n12915), .A2(n12914), .ZN(n4712) );
  OAI22_X2 U14990 ( .A1(n13363), .A2(n12916), .B1(n5583), .B2(n13430), .ZN(
        n4715) );
  INV_X4 U14991 ( .A(n12918), .ZN(n12920) );
  NAND2_X2 U14992 ( .A1(n6581), .A2(ifInst[26]), .ZN(n13428) );
  NAND2_X2 U14993 ( .A1(n6587), .A2(idOut_16_), .ZN(n12919) );
  INV_X4 U14994 ( .A(ifInst[31]), .ZN(n13497) );
  NAND2_X2 U14995 ( .A1(n13430), .A2(n13363), .ZN(n13399) );
  NAND2_X2 U14996 ( .A1(n13399), .A2(n13430), .ZN(n13332) );
  NAND2_X2 U14997 ( .A1(n6587), .A2(idOut_28_), .ZN(n12922) );
  INV_X4 U14998 ( .A(n12924), .ZN(n12930) );
  NAND2_X2 U14999 ( .A1(n5306), .A2(daddr[20]), .ZN(n12929) );
  NAND2_X2 U15000 ( .A1(dwData[20]), .A2(n6609), .ZN(n12928) );
  OAI211_X2 U15001 ( .C1(n12930), .C2(n6578), .A(n12929), .B(n12928), .ZN(
        n13646) );
  INV_X4 U15002 ( .A(n12931), .ZN(n12934) );
  NAND2_X2 U15003 ( .A1(n5306), .A2(daddr[19]), .ZN(n12933) );
  NAND2_X2 U15004 ( .A1(dwData[19]), .A2(n6609), .ZN(n12932) );
  OAI211_X2 U15005 ( .C1(n12934), .C2(n6578), .A(n12933), .B(n12932), .ZN(
        n13645) );
  INV_X4 U15006 ( .A(n12935), .ZN(n12938) );
  NAND2_X2 U15007 ( .A1(n5306), .A2(daddr[15]), .ZN(n12937) );
  NAND2_X2 U15008 ( .A1(dwData[15]), .A2(n6610), .ZN(n12936) );
  OAI211_X2 U15009 ( .C1(n12938), .C2(n6578), .A(n12937), .B(n12936), .ZN(
        n13641) );
  NOR2_X4 U15010 ( .A1(n12941), .A2(n6555), .ZN(n12942) );
  NOR3_X4 U15011 ( .A1(n5035), .A2(n12943), .A3(n12942), .ZN(n12949) );
  NAND2_X2 U15012 ( .A1(aluBoi_aluBoi_shft_sraout[15]), .A2(n5460), .ZN(n12948) );
  AOI22_X2 U15013 ( .A1(n12946), .A2(n13062), .B1(aluBoi_multBoi_temppp[12]), 
        .B2(net368069), .ZN(n12947) );
  INV_X4 U15014 ( .A(n12950), .ZN(n12953) );
  NAND2_X2 U15015 ( .A1(n5306), .A2(daddr[14]), .ZN(n12952) );
  NAND2_X2 U15016 ( .A1(dwData[14]), .A2(n6610), .ZN(n12951) );
  OAI211_X2 U15017 ( .C1(n12953), .C2(n6578), .A(n12952), .B(n12951), .ZN(
        n13640) );
  INV_X4 U15018 ( .A(n12954), .ZN(n12957) );
  NAND2_X2 U15019 ( .A1(n5306), .A2(daddr[10]), .ZN(n12956) );
  NAND2_X2 U15020 ( .A1(dwData[10]), .A2(n6610), .ZN(n12955) );
  OAI211_X2 U15021 ( .C1(n12957), .C2(n6578), .A(n12956), .B(n12955), .ZN(
        n13636) );
  INV_X4 U15022 ( .A(n12958), .ZN(n12959) );
  AOI22_X2 U15023 ( .A1(n13019), .A2(n12959), .B1(aluBoi_multBoi_temppp[7]), 
        .B2(net368069), .ZN(n12964) );
  NAND2_X2 U15024 ( .A1(aluBoi_aluBoi_shft_sraout[10]), .A2(n5460), .ZN(n12963) );
  NAND2_X2 U15025 ( .A1(daddr[10]), .A2(n6610), .ZN(n12962) );
  AOI22_X2 U15026 ( .A1(n13062), .A2(n12960), .B1(
        aluBoi_aluBoi_shft_sllout[10]), .B2(n5315), .ZN(n12961) );
  NAND4_X2 U15027 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n4726) );
  INV_X4 U15028 ( .A(n12965), .ZN(n12968) );
  NAND2_X2 U15029 ( .A1(n5306), .A2(daddr[9]), .ZN(n12967) );
  NAND2_X2 U15030 ( .A1(dwData[9]), .A2(n6610), .ZN(n12966) );
  OAI211_X2 U15031 ( .C1(n12968), .C2(n6578), .A(n12967), .B(n12966), .ZN(
        n13635) );
  NAND2_X2 U15032 ( .A1(n5306), .A2(daddr[5]), .ZN(n12971) );
  NAND2_X2 U15033 ( .A1(dwData[5]), .A2(n6610), .ZN(n12970) );
  OAI211_X2 U15034 ( .C1(n12972), .C2(n6578), .A(n12971), .B(n12970), .ZN(
        n13631) );
  INV_X4 U15035 ( .A(n12973), .ZN(n12974) );
  AOI22_X2 U15036 ( .A1(n13019), .A2(n12974), .B1(aluBoi_multBoi_temppp[2]), 
        .B2(net368069), .ZN(n12979) );
  NAND2_X2 U15037 ( .A1(aluBoi_aluBoi_shft_sraout[5]), .A2(n5460), .ZN(n12978)
         );
  NAND2_X2 U15038 ( .A1(daddr[5]), .A2(n6610), .ZN(n12977) );
  AOI22_X2 U15039 ( .A1(aluBoi_aluBoi_shft_sllout[5]), .A2(n5315), .B1(n6605), 
        .B2(n12975), .ZN(n12976) );
  NAND4_X2 U15040 ( .A1(n12979), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n4729) );
  INV_X4 U15041 ( .A(n13514), .ZN(n12982) );
  INV_X4 U15042 ( .A(n12980), .ZN(n12981) );
  AOI22_X2 U15043 ( .A1(n12982), .A2(n12981), .B1(aluBoi_multBoi_temppp[6]), 
        .B2(net368069), .ZN(n12987) );
  NAND2_X2 U15044 ( .A1(aluBoi_aluBoi_shft_sraout[9]), .A2(n5460), .ZN(n12986)
         );
  NAND2_X2 U15045 ( .A1(daddr[9]), .A2(n6610), .ZN(n12985) );
  AOI22_X2 U15046 ( .A1(n13062), .A2(n12983), .B1(aluBoi_aluBoi_shft_sllout[9]), .B2(n5315), .ZN(n12984) );
  NAND4_X2 U15047 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        n4730) );
  INV_X4 U15048 ( .A(n12988), .ZN(n12991) );
  NAND2_X2 U15049 ( .A1(n5306), .A2(daddr[8]), .ZN(n12990) );
  NAND2_X2 U15050 ( .A1(dwData[8]), .A2(n6610), .ZN(n12989) );
  OAI211_X2 U15051 ( .C1(n12991), .C2(n6578), .A(n12990), .B(n12989), .ZN(
        n13634) );
  MUX2_X2 U15052 ( .A(n12993), .B(n12992), .S(n6821), .Z(n12997) );
  MUX2_X2 U15053 ( .A(n12995), .B(n12994), .S(n6821), .Z(n12996) );
  MUX2_X2 U15054 ( .A(n12997), .B(n12996), .S(n6830), .Z(n13005) );
  MUX2_X2 U15055 ( .A(n12999), .B(n12998), .S(n6821), .Z(n13003) );
  MUX2_X2 U15056 ( .A(n13001), .B(n13000), .S(n6821), .Z(n13002) );
  MUX2_X2 U15057 ( .A(n13003), .B(n13002), .S(n6830), .Z(n13004) );
  MUX2_X2 U15058 ( .A(n13005), .B(n13004), .S(n6834), .Z(n13006) );
  INV_X4 U15059 ( .A(n13006), .ZN(n13009) );
  NAND2_X2 U15060 ( .A1(n5306), .A2(daddr[4]), .ZN(n13008) );
  NAND2_X2 U15061 ( .A1(dwData[4]), .A2(n6610), .ZN(n13007) );
  OAI211_X2 U15062 ( .C1(n13009), .C2(n6578), .A(n13008), .B(n13007), .ZN(
        n13630) );
  INV_X4 U15063 ( .A(n13010), .ZN(n13011) );
  AOI22_X2 U15064 ( .A1(n13019), .A2(n13011), .B1(aluBoi_multBoi_temppp[1]), 
        .B2(net368069), .ZN(n13016) );
  NAND2_X2 U15065 ( .A1(aluBoi_aluBoi_shft_sraout[4]), .A2(n5460), .ZN(n13015)
         );
  AOI22_X2 U15066 ( .A1(daddr[4]), .A2(n6609), .B1(
        aluBoi_aluBoi_shft_sllout[4]), .B2(n5315), .ZN(n13014) );
  NAND2_X2 U15067 ( .A1(n6605), .A2(n13012), .ZN(n13013) );
  NAND4_X2 U15068 ( .A1(n13016), .A2(n13015), .A3(n13014), .A4(n13013), .ZN(
        n4733) );
  INV_X4 U15069 ( .A(n6555), .ZN(n13019) );
  INV_X4 U15070 ( .A(n13017), .ZN(n13018) );
  AOI22_X2 U15071 ( .A1(n13019), .A2(n13018), .B1(aluBoi_multBoi_temppp[5]), 
        .B2(net368069), .ZN(n13024) );
  NAND2_X2 U15072 ( .A1(aluBoi_aluBoi_shft_sraout[8]), .A2(n5460), .ZN(n13023)
         );
  NAND2_X2 U15073 ( .A1(daddr[8]), .A2(n6610), .ZN(n13022) );
  AOI22_X2 U15074 ( .A1(n13062), .A2(n13020), .B1(aluBoi_aluBoi_shft_sllout[8]), .B2(n5315), .ZN(n13021) );
  NAND4_X2 U15075 ( .A1(n13024), .A2(n13023), .A3(n13022), .A4(n13021), .ZN(
        n4734) );
  INV_X4 U15076 ( .A(n13025), .ZN(n13028) );
  NAND2_X2 U15077 ( .A1(n5306), .A2(daddr[7]), .ZN(n13027) );
  NAND2_X2 U15078 ( .A1(dwData[7]), .A2(n6610), .ZN(n13026) );
  OAI211_X2 U15079 ( .C1(n13028), .C2(n6578), .A(n13027), .B(n13026), .ZN(
        n13633) );
  INV_X4 U15080 ( .A(n13029), .ZN(n13030) );
  AOI22_X2 U15081 ( .A1(n12982), .A2(n13030), .B1(aluBoi_multBoi_temppp[4]), 
        .B2(net368069), .ZN(n13035) );
  NAND2_X2 U15082 ( .A1(aluBoi_aluBoi_shft_sraout[7]), .A2(n5460), .ZN(n13034)
         );
  NAND2_X2 U15083 ( .A1(daddr[7]), .A2(n6610), .ZN(n13033) );
  AOI22_X2 U15084 ( .A1(n13062), .A2(n13031), .B1(aluBoi_aluBoi_shft_sllout[7]), .B2(n5315), .ZN(n13032) );
  NAND4_X2 U15085 ( .A1(n13035), .A2(n13034), .A3(n13033), .A4(n13032), .ZN(
        n4736) );
  NAND2_X2 U15086 ( .A1(n5306), .A2(daddr[6]), .ZN(n13038) );
  NAND2_X2 U15087 ( .A1(dwData[6]), .A2(n6610), .ZN(n13037) );
  OAI211_X2 U15088 ( .C1(n13039), .C2(n6578), .A(n13038), .B(n13037), .ZN(
        n13632) );
  INV_X4 U15089 ( .A(n13040), .ZN(n13041) );
  AOI22_X2 U15090 ( .A1(n12982), .A2(n13041), .B1(aluBoi_multBoi_temppp[3]), 
        .B2(net368069), .ZN(n13046) );
  NAND2_X2 U15091 ( .A1(aluBoi_aluBoi_shft_sraout[6]), .A2(n5460), .ZN(n13045)
         );
  NAND2_X2 U15092 ( .A1(daddr[6]), .A2(n6610), .ZN(n13044) );
  AOI22_X2 U15093 ( .A1(aluBoi_aluBoi_shft_sllout[6]), .A2(n5315), .B1(n6605), 
        .B2(n13042), .ZN(n13043) );
  NAND4_X2 U15094 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n4738) );
  INV_X4 U15095 ( .A(n13047), .ZN(n13048) );
  AOI22_X2 U15096 ( .A1(n12982), .A2(n13048), .B1(aluBoi_multBoi_temppp[11]), 
        .B2(net368069), .ZN(n13054) );
  NAND2_X2 U15097 ( .A1(aluBoi_aluBoi_shft_sraout[14]), .A2(n5460), .ZN(n13053) );
  NAND2_X2 U15098 ( .A1(daddr[14]), .A2(n6610), .ZN(n13052) );
  AOI22_X2 U15099 ( .A1(n13062), .A2(n13050), .B1(
        aluBoi_aluBoi_shft_sllout[14]), .B2(n5315), .ZN(n13051) );
  NAND4_X2 U15100 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n4739) );
  INV_X4 U15101 ( .A(n13055), .ZN(n13058) );
  NAND2_X2 U15102 ( .A1(n5306), .A2(daddr[13]), .ZN(n13057) );
  NAND2_X2 U15103 ( .A1(dwData[13]), .A2(n6610), .ZN(n13056) );
  OAI211_X2 U15104 ( .C1(n13058), .C2(n6578), .A(n13057), .B(n13056), .ZN(
        n13639) );
  INV_X4 U15105 ( .A(n13059), .ZN(n13060) );
  AOI22_X2 U15106 ( .A1(n12982), .A2(n13060), .B1(aluBoi_multBoi_temppp[10]), 
        .B2(net368069), .ZN(n13066) );
  NAND2_X2 U15107 ( .A1(aluBoi_aluBoi_shft_sraout[13]), .A2(n5460), .ZN(n13065) );
  NAND2_X2 U15108 ( .A1(daddr[13]), .A2(n6610), .ZN(n13064) );
  AOI22_X2 U15109 ( .A1(n13062), .A2(n13061), .B1(
        aluBoi_aluBoi_shft_sllout[13]), .B2(n5315), .ZN(n13063) );
  NAND4_X2 U15110 ( .A1(n13066), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        n4741) );
  INV_X4 U15111 ( .A(n13067), .ZN(n13070) );
  NAND2_X2 U15112 ( .A1(n5306), .A2(daddr[12]), .ZN(n13069) );
  NAND2_X2 U15113 ( .A1(dwData[12]), .A2(n6610), .ZN(n13068) );
  OAI211_X2 U15114 ( .C1(n13070), .C2(n6578), .A(n13069), .B(n13068), .ZN(
        n13638) );
  INV_X4 U15115 ( .A(n13071), .ZN(n13072) );
  AOI22_X2 U15116 ( .A1(n13019), .A2(n13072), .B1(aluBoi_multBoi_temppp[9]), 
        .B2(net368069), .ZN(n13078) );
  NAND2_X2 U15117 ( .A1(aluBoi_aluBoi_shft_sraout[12]), .A2(n5460), .ZN(n13077) );
  NAND2_X2 U15118 ( .A1(daddr[12]), .A2(n6610), .ZN(n13076) );
  INV_X4 U15119 ( .A(n13073), .ZN(n13074) );
  AOI22_X2 U15120 ( .A1(n13062), .A2(n13074), .B1(
        aluBoi_aluBoi_shft_sllout[12]), .B2(n5315), .ZN(n13075) );
  NAND4_X2 U15121 ( .A1(n13078), .A2(n13077), .A3(n13076), .A4(n13075), .ZN(
        n4743) );
  INV_X4 U15122 ( .A(n13079), .ZN(n13082) );
  NAND2_X2 U15123 ( .A1(n5306), .A2(daddr[11]), .ZN(n13081) );
  NAND2_X2 U15124 ( .A1(dwData[11]), .A2(n6610), .ZN(n13080) );
  OAI211_X2 U15125 ( .C1(n13082), .C2(n6578), .A(n13081), .B(n13080), .ZN(
        n13637) );
  INV_X4 U15126 ( .A(n13083), .ZN(n13084) );
  AOI22_X2 U15127 ( .A1(n13019), .A2(n13084), .B1(aluBoi_multBoi_temppp[8]), 
        .B2(net368069), .ZN(n13089) );
  NAND2_X2 U15128 ( .A1(aluBoi_aluBoi_shft_sraout[11]), .A2(n5460), .ZN(n13088) );
  NAND2_X2 U15129 ( .A1(daddr[11]), .A2(n6610), .ZN(n13087) );
  AOI22_X2 U15130 ( .A1(n6605), .A2(n13085), .B1(aluBoi_aluBoi_shft_sllout[11]), .B2(n5315), .ZN(n13086) );
  NAND4_X2 U15131 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n4745) );
  INV_X4 U15132 ( .A(n13090), .ZN(n13091) );
  NAND2_X2 U15133 ( .A1(aluBoi_aluBoi_shft_sraout[19]), .A2(n5460), .ZN(n13095) );
  NAND2_X2 U15134 ( .A1(daddr[19]), .A2(n6610), .ZN(n13094) );
  AOI22_X2 U15135 ( .A1(n6605), .A2(n13092), .B1(aluBoi_aluBoi_shft_sllout[19]), .B2(n5315), .ZN(n13093) );
  NAND4_X2 U15136 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        n4746) );
  INV_X4 U15137 ( .A(n13097), .ZN(n13100) );
  NAND2_X2 U15138 ( .A1(n5306), .A2(daddr[18]), .ZN(n13099) );
  NAND2_X2 U15139 ( .A1(dwData[18]), .A2(n6610), .ZN(n13098) );
  OAI211_X2 U15140 ( .C1(n13100), .C2(n6578), .A(n13099), .B(n13098), .ZN(
        n13644) );
  AOI222_X4 U15141 ( .A1(n12982), .A2(n9063), .B1(aluBoi_multBoi_temppp[15]), 
        .B2(net368069), .C1(n5316), .C2(n6074), .ZN(n13106) );
  NAND2_X2 U15142 ( .A1(aluBoi_aluBoi_shft_sraout[18]), .A2(n5460), .ZN(n13105) );
  NAND2_X2 U15143 ( .A1(daddr[18]), .A2(n6610), .ZN(n13104) );
  AOI22_X2 U15144 ( .A1(n6605), .A2(n13102), .B1(aluBoi_aluBoi_shft_sllout[18]), .B2(n5315), .ZN(n13103) );
  NAND4_X2 U15145 ( .A1(n13106), .A2(n13105), .A3(n13104), .A4(n13103), .ZN(
        n4748) );
  INV_X4 U15146 ( .A(n13107), .ZN(n13110) );
  NAND2_X2 U15147 ( .A1(n5306), .A2(daddr[17]), .ZN(n13109) );
  NAND2_X2 U15148 ( .A1(dwData[17]), .A2(n6610), .ZN(n13108) );
  OAI211_X2 U15149 ( .C1(n13110), .C2(n6578), .A(n13109), .B(n13108), .ZN(
        n13643) );
  INV_X4 U15150 ( .A(n13111), .ZN(n13112) );
  NAND2_X2 U15151 ( .A1(aluBoi_aluBoi_shft_sraout[17]), .A2(n5460), .ZN(n13116) );
  NAND2_X2 U15152 ( .A1(daddr[17]), .A2(n6610), .ZN(n13115) );
  AOI22_X2 U15153 ( .A1(n6605), .A2(n13113), .B1(aluBoi_aluBoi_shft_sllout[17]), .B2(n5315), .ZN(n13114) );
  NAND4_X2 U15154 ( .A1(n13117), .A2(n13116), .A3(n13115), .A4(n13114), .ZN(
        n4750) );
  INV_X4 U15155 ( .A(n13118), .ZN(n13121) );
  NAND2_X2 U15156 ( .A1(n5306), .A2(daddr[16]), .ZN(n13120) );
  NAND2_X2 U15157 ( .A1(dwData[16]), .A2(n6610), .ZN(n13119) );
  OAI211_X2 U15158 ( .C1(n13121), .C2(n6578), .A(n13120), .B(n13119), .ZN(
        n13642) );
  INV_X4 U15159 ( .A(n13122), .ZN(n13123) );
  NAND2_X2 U15160 ( .A1(aluBoi_aluBoi_shft_sraout[16]), .A2(n5460), .ZN(n13127) );
  NAND2_X2 U15161 ( .A1(daddr[16]), .A2(n6610), .ZN(n13126) );
  AOI22_X2 U15162 ( .A1(n6605), .A2(n13124), .B1(aluBoi_aluBoi_shft_sllout[16]), .B2(n5315), .ZN(n13125) );
  NAND4_X2 U15163 ( .A1(n13128), .A2(n13127), .A3(n13126), .A4(n13125), .ZN(
        n4752) );
  INV_X4 U15164 ( .A(n13129), .ZN(n13130) );
  NAND2_X2 U15165 ( .A1(aluBoi_aluBoi_shft_sraout[20]), .A2(n5460), .ZN(n13134) );
  NAND2_X2 U15166 ( .A1(daddr[20]), .A2(n6610), .ZN(n13133) );
  AOI22_X2 U15167 ( .A1(n6605), .A2(n13131), .B1(aluBoi_aluBoi_shft_sllout[20]), .B2(n5315), .ZN(n13132) );
  NAND4_X2 U15168 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n4753) );
  INV_X4 U15169 ( .A(n13136), .ZN(n13139) );
  NAND2_X2 U15170 ( .A1(n5306), .A2(daddr[21]), .ZN(n13138) );
  NAND2_X2 U15171 ( .A1(dwData[21]), .A2(n6610), .ZN(n13137) );
  OAI211_X2 U15172 ( .C1(n13139), .C2(n6578), .A(n13138), .B(n13137), .ZN(
        n13647) );
  NAND2_X2 U15173 ( .A1(aluBoi_aluBoi_shft_sraout[21]), .A2(n5460), .ZN(n13145) );
  NAND2_X2 U15174 ( .A1(daddr[21]), .A2(n6610), .ZN(n13144) );
  AOI22_X2 U15175 ( .A1(n6605), .A2(n13142), .B1(aluBoi_aluBoi_shft_sllout[21]), .B2(n5315), .ZN(n13143) );
  NAND4_X2 U15176 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        n4755) );
  INV_X4 U15177 ( .A(n13147), .ZN(n13150) );
  NAND2_X2 U15178 ( .A1(n5306), .A2(daddr[22]), .ZN(n13149) );
  NAND2_X2 U15179 ( .A1(dwData[22]), .A2(n6610), .ZN(n13148) );
  OAI211_X2 U15180 ( .C1(n13150), .C2(n6578), .A(n13149), .B(n13148), .ZN(
        n13648) );
  NAND2_X2 U15181 ( .A1(aluBoi_multBoi_temppp[19]), .A2(net368069), .ZN(n13156) );
  NAND2_X2 U15182 ( .A1(daddr[22]), .A2(n6609), .ZN(n13155) );
  NAND2_X2 U15183 ( .A1(n5316), .A2(aluBoi_imm32w_6_), .ZN(n13153) );
  NAND4_X2 U15184 ( .A1(n13154), .A2(n13155), .A3(n13156), .A4(n13153), .ZN(
        n4757) );
  INV_X4 U15185 ( .A(n13157), .ZN(n13160) );
  NAND2_X2 U15186 ( .A1(n5306), .A2(daddr[23]), .ZN(n13159) );
  NAND2_X2 U15187 ( .A1(dwData[23]), .A2(n6610), .ZN(n13158) );
  OAI211_X2 U15188 ( .C1(n13160), .C2(n6578), .A(n13159), .B(n13158), .ZN(
        n13649) );
  NAND2_X2 U15189 ( .A1(aluBoi_multBoi_temppp[20]), .A2(net368069), .ZN(n13166) );
  NAND2_X2 U15190 ( .A1(daddr[23]), .A2(n6609), .ZN(n13165) );
  NAND2_X2 U15191 ( .A1(n5316), .A2(aluBoi_imm32w_7_), .ZN(n13163) );
  NAND4_X2 U15192 ( .A1(n13166), .A2(n13165), .A3(n13164), .A4(n13163), .ZN(
        n4759) );
  INV_X4 U15193 ( .A(n13167), .ZN(n13170) );
  NAND2_X2 U15194 ( .A1(n5306), .A2(daddr[25]), .ZN(n13169) );
  NAND2_X2 U15195 ( .A1(dwData[25]), .A2(n6610), .ZN(n13168) );
  OAI211_X2 U15196 ( .C1(n13170), .C2(n6578), .A(n13169), .B(n13168), .ZN(
        n13651) );
  NAND2_X2 U15197 ( .A1(aluBoi_multBoi_temppp[22]), .A2(net368069), .ZN(n13176) );
  NAND2_X2 U15198 ( .A1(daddr[25]), .A2(n6609), .ZN(n13175) );
  OAI21_X4 U15199 ( .B1(n13172), .B2(n13171), .A(n13062), .ZN(n13174) );
  NAND2_X2 U15200 ( .A1(n5316), .A2(aluBoi_imm32w_9_), .ZN(n13173) );
  NAND4_X2 U15201 ( .A1(n13174), .A2(n13175), .A3(n13176), .A4(n13173), .ZN(
        n4761) );
  INV_X4 U15202 ( .A(n13177), .ZN(n13180) );
  NAND2_X2 U15203 ( .A1(n5306), .A2(daddr[24]), .ZN(n13179) );
  NAND2_X2 U15204 ( .A1(dwData[24]), .A2(n6610), .ZN(n13178) );
  OAI211_X2 U15205 ( .C1(n13180), .C2(n13375), .A(n13179), .B(n13178), .ZN(
        n13650) );
  NAND2_X2 U15206 ( .A1(aluBoi_multBoi_temppp[21]), .A2(net368069), .ZN(n13186) );
  NAND2_X2 U15207 ( .A1(daddr[24]), .A2(n6609), .ZN(n13185) );
  NAND2_X2 U15208 ( .A1(n5316), .A2(aluBoi_imm32w_8_), .ZN(n13183) );
  NAND4_X2 U15209 ( .A1(n13186), .A2(n13185), .A3(n13184), .A4(n13183), .ZN(
        n4763) );
  INV_X4 U15210 ( .A(n13187), .ZN(n13190) );
  NAND2_X2 U15211 ( .A1(n5306), .A2(daddr[28]), .ZN(n13189) );
  NAND2_X2 U15212 ( .A1(dwData[28]), .A2(n6610), .ZN(n13188) );
  OAI211_X2 U15213 ( .C1(n13190), .C2(n13375), .A(n13189), .B(n13188), .ZN(
        n13654) );
  NOR2_X4 U15214 ( .A1(n13192), .A2(n13191), .ZN(n13194) );
  INV_X4 U15215 ( .A(n13195), .ZN(n13198) );
  NAND2_X2 U15216 ( .A1(n5306), .A2(daddr[27]), .ZN(n13197) );
  NAND2_X2 U15217 ( .A1(dwData[27]), .A2(n6610), .ZN(n13196) );
  OAI211_X2 U15218 ( .C1(n13198), .C2(n13375), .A(n13197), .B(n13196), .ZN(
        n13653) );
  NAND2_X2 U15219 ( .A1(aluBoi_multBoi_temppp[24]), .A2(net368069), .ZN(n13204) );
  NAND2_X2 U15220 ( .A1(daddr[27]), .A2(n6609), .ZN(n13203) );
  NAND2_X2 U15221 ( .A1(n5316), .A2(aluBoi_imm32w_11_), .ZN(n13201) );
  NAND4_X2 U15222 ( .A1(n13202), .A2(n13203), .A3(n13204), .A4(n13201), .ZN(
        n4767) );
  INV_X4 U15223 ( .A(n13205), .ZN(n13208) );
  NAND2_X2 U15224 ( .A1(n5306), .A2(daddr[26]), .ZN(n13207) );
  NAND2_X2 U15225 ( .A1(dwData[26]), .A2(n6609), .ZN(n13206) );
  OAI211_X2 U15226 ( .C1(n13208), .C2(n13375), .A(n13207), .B(n13206), .ZN(
        n13652) );
  NAND2_X2 U15227 ( .A1(aluBoi_multBoi_temppp[23]), .A2(net368069), .ZN(n13214) );
  NAND2_X2 U15228 ( .A1(daddr[26]), .A2(n6609), .ZN(n13213) );
  NAND2_X2 U15229 ( .A1(n5316), .A2(aluBoi_imm32w_10_), .ZN(n13211) );
  NAND4_X2 U15230 ( .A1(n13214), .A2(n13213), .A3(n13212), .A4(n13211), .ZN(
        n4769) );
  INV_X4 U15231 ( .A(n13215), .ZN(n13218) );
  NAND2_X2 U15232 ( .A1(n5306), .A2(daddr[30]), .ZN(n13217) );
  NAND2_X2 U15233 ( .A1(dwData[30]), .A2(n6609), .ZN(n13216) );
  OAI211_X2 U15234 ( .C1(n13218), .C2(n13375), .A(n13217), .B(n13216), .ZN(
        n13656) );
  INV_X4 U15235 ( .A(n13219), .ZN(n13221) );
  INV_X4 U15236 ( .A(n13223), .ZN(n13225) );
  NOR2_X4 U15237 ( .A1(n13225), .A2(n13224), .ZN(n13227) );
  NAND2_X2 U15238 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  INV_X4 U15239 ( .A(n13233), .ZN(n13236) );
  NAND2_X2 U15240 ( .A1(n5306), .A2(daddr[29]), .ZN(n13235) );
  NAND2_X2 U15241 ( .A1(dwData[29]), .A2(n6609), .ZN(n13234) );
  OAI211_X2 U15242 ( .C1(n13236), .C2(n13375), .A(n13235), .B(n13234), .ZN(
        n13655) );
  NAND2_X2 U15243 ( .A1(n5316), .A2(aluBoi_imm32w_13_), .ZN(n13242) );
  NAND2_X2 U15244 ( .A1(aluBoi_multBoi_temppp[26]), .A2(net368069), .ZN(n13240) );
  NAND2_X2 U15245 ( .A1(daddr[29]), .A2(n6609), .ZN(n13239) );
  NAND4_X2 U15246 ( .A1(n13241), .A2(n13242), .A3(n13240), .A4(n13239), .ZN(
        n4773) );
  NAND2_X2 U15247 ( .A1(n5306), .A2(daddr[3]), .ZN(n13245) );
  NAND2_X2 U15248 ( .A1(dwData[3]), .A2(n6609), .ZN(n13244) );
  OAI211_X2 U15249 ( .C1(n13246), .C2(n13375), .A(n13245), .B(n13244), .ZN(
        n13629) );
  INV_X4 U15250 ( .A(n13247), .ZN(n13248) );
  NOR2_X4 U15251 ( .A1(n6554), .A2(n13248), .ZN(n13249) );
  NAND2_X2 U15252 ( .A1(aluBoi_aluBoi_shft_sraout[3]), .A2(n5460), .ZN(n13253)
         );
  NAND2_X2 U15253 ( .A1(daddr[3]), .A2(n6609), .ZN(n13252) );
  AOI22_X2 U15254 ( .A1(n6605), .A2(n13250), .B1(aluBoi_aluBoi_shft_sllout[3]), 
        .B2(n5315), .ZN(n13251) );
  NAND4_X2 U15255 ( .A1(n13254), .A2(n13253), .A3(n13252), .A4(n13251), .ZN(
        n4775) );
  NAND2_X2 U15256 ( .A1(n5306), .A2(daddr[2]), .ZN(n13257) );
  NAND2_X2 U15257 ( .A1(dwData[2]), .A2(n6609), .ZN(n13256) );
  OAI211_X2 U15258 ( .C1(n13258), .C2(n13375), .A(n13257), .B(n13256), .ZN(
        n13660) );
  NAND2_X2 U15259 ( .A1(n6605), .A2(n13259), .ZN(n13265) );
  NAND2_X2 U15260 ( .A1(aluBoi_aluBoi_shft_sllout[2]), .A2(n5315), .ZN(n13264)
         );
  NAND2_X2 U15261 ( .A1(daddr[2]), .A2(n6609), .ZN(n13263) );
  NOR2_X4 U15262 ( .A1(n13260), .A2(n13514), .ZN(n13261) );
  NAND4_X2 U15263 ( .A1(n13265), .A2(n13264), .A3(n13263), .A4(n13262), .ZN(
        n4777) );
  INV_X4 U15264 ( .A(n13266), .ZN(n13269) );
  NAND2_X2 U15265 ( .A1(n5306), .A2(daddr[1]), .ZN(n13268) );
  NAND2_X2 U15266 ( .A1(dwData[1]), .A2(n6609), .ZN(n13267) );
  NAND2_X2 U15267 ( .A1(n6605), .A2(n13270), .ZN(n13276) );
  NAND2_X2 U15268 ( .A1(aluBoi_aluBoi_shft_sllout[1]), .A2(n5315), .ZN(n13275)
         );
  NAND2_X2 U15269 ( .A1(daddr[1]), .A2(n6609), .ZN(n13274) );
  NOR2_X4 U15270 ( .A1(n13271), .A2(n6554), .ZN(n13272) );
  NAND4_X2 U15271 ( .A1(n13276), .A2(n13275), .A3(n13274), .A4(n13273), .ZN(
        n4779) );
  INV_X4 U15272 ( .A(n13277), .ZN(n13280) );
  NAND2_X2 U15273 ( .A1(n5306), .A2(daddr[0]), .ZN(n13279) );
  NAND2_X2 U15274 ( .A1(dwData[0]), .A2(n6609), .ZN(n13278) );
  OAI211_X2 U15275 ( .C1(n13280), .C2(n13375), .A(n13279), .B(n13278), .ZN(
        n13658) );
  NAND2_X2 U15276 ( .A1(aluBoi_aluBoi_shft_sraout[0]), .A2(n5460), .ZN(n13287)
         );
  INV_X4 U15277 ( .A(aluBoi_condOut_0_), .ZN(n13281) );
  AOI21_X4 U15278 ( .B1(n13282), .B2(n6608), .A(net358577), .ZN(n13286) );
  NAND2_X2 U15279 ( .A1(daddr[0]), .A2(n6609), .ZN(n13285) );
  AOI22_X2 U15280 ( .A1(n13062), .A2(n13283), .B1(aluBoi_aluBoi_shft_sllout[0]), .B2(n5315), .ZN(n13284) );
  NAND4_X2 U15281 ( .A1(n13287), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n4781) );
  INV_X4 U15282 ( .A(n13308), .ZN(n13289) );
  INV_X4 U15283 ( .A(ifInst[1]), .ZN(n13499) );
  MUX2_X2 U15284 ( .A(n13499), .B(n13302), .S(ifInst[2]), .Z(n13290) );
  INV_X4 U15285 ( .A(n13400), .ZN(n13295) );
  NAND2_X2 U15286 ( .A1(n6581), .A2(n13294), .ZN(n13299) );
  NAND2_X2 U15287 ( .A1(n6581), .A2(n13493), .ZN(n13434) );
  INV_X4 U15288 ( .A(n13434), .ZN(n13296) );
  NAND3_X4 U15289 ( .A1(n13296), .A2(ifInst[27]), .A3(n13295), .ZN(n13298) );
  NAND2_X2 U15290 ( .A1(idOut_21_), .A2(n6588), .ZN(n13297) );
  INV_X4 U15291 ( .A(n2054), .ZN(n13300) );
  AOI22_X2 U15292 ( .A1(n13302), .A2(n13289), .B1(n13301), .B2(n13300), .ZN(
        n13305) );
  INV_X4 U15293 ( .A(n13428), .ZN(n13351) );
  NAND4_X2 U15294 ( .A1(ifInst[28]), .A2(ifInst[30]), .A3(n13351), .A4(n13321), 
        .ZN(n13311) );
  NAND2_X2 U15295 ( .A1(n5492), .A2(idOut_24_), .ZN(n13304) );
  OAI211_X2 U15296 ( .C1(n13305), .C2(n13363), .A(n13311), .B(n13304), .ZN(
        n4783) );
  NAND2_X2 U15297 ( .A1(ifInst[27]), .A2(n13539), .ZN(n13325) );
  INV_X4 U15298 ( .A(n13325), .ZN(n13306) );
  NAND2_X2 U15299 ( .A1(n5380), .A2(n6582), .ZN(n13425) );
  NAND2_X2 U15300 ( .A1(n13306), .A2(n13365), .ZN(n13312) );
  NAND2_X2 U15301 ( .A1(n13307), .A2(n5343), .ZN(n13366) );
  MUX2_X2 U15302 ( .A(n13366), .B(n13308), .S(ifInst[0]), .Z(n13309) );
  NAND2_X2 U15303 ( .A1(n6581), .A2(ifInst[1]), .ZN(n13408) );
  NAND2_X2 U15304 ( .A1(n6587), .A2(idOut_22_), .ZN(n13310) );
  NAND4_X2 U15305 ( .A1(n13312), .A2(n5700), .A3(n13311), .A4(n13310), .ZN(
        n4784) );
  INV_X4 U15306 ( .A(n13433), .ZN(n13396) );
  NAND2_X2 U15307 ( .A1(n13314), .A2(n13313), .ZN(n13316) );
  NAND2_X2 U15308 ( .A1(n2013), .A2(n2011), .ZN(n13315) );
  NOR4_X2 U15309 ( .A1(n13316), .A2(n13315), .A3(n2009), .A4(n5561), .ZN(
        n13318) );
  MUX2_X2 U15310 ( .A(n13318), .B(n13317), .S(ifInst[0]), .Z(n13320) );
  NAND4_X2 U15311 ( .A1(n13396), .A2(n13320), .A3(n5346), .A4(n13319), .ZN(
        n13329) );
  INV_X4 U15312 ( .A(n13322), .ZN(n13323) );
  NAND2_X2 U15313 ( .A1(n13323), .A2(n13497), .ZN(n13429) );
  INV_X4 U15314 ( .A(n13429), .ZN(n13326) );
  INV_X4 U15315 ( .A(n13324), .ZN(n13422) );
  NAND4_X2 U15316 ( .A1(n13329), .A2(n13399), .A3(n13328), .A4(n13327), .ZN(
        n13331) );
  NAND2_X2 U15317 ( .A1(idRegWr), .A2(n6588), .ZN(n13330) );
  NAND2_X2 U15318 ( .A1(n13331), .A2(n13330), .ZN(n4786) );
  OAI22_X2 U15319 ( .A1(n5714), .A2(n13430), .B1(n13333), .B2(n13332), .ZN(
        n4787) );
  NAND2_X2 U15320 ( .A1(n13334), .A2(n5312), .ZN(n13357) );
  INV_X4 U15321 ( .A(n13335), .ZN(n13336) );
  NAND2_X2 U15322 ( .A1(n13360), .A2(n13336), .ZN(n13338) );
  NAND2_X2 U15323 ( .A1(idOut_18_), .A2(n6589), .ZN(n13337) );
  OAI211_X2 U15324 ( .C1(n13357), .C2(n13339), .A(n13338), .B(n13337), .ZN(
        n4788) );
  INV_X4 U15325 ( .A(n13340), .ZN(n13342) );
  INV_X4 U15326 ( .A(n13348), .ZN(n13343) );
  OAI21_X4 U15327 ( .B1(n13345), .B2(n13344), .A(n6581), .ZN(n13347) );
  NAND2_X2 U15328 ( .A1(n6587), .A2(idOut_19_), .ZN(n13346) );
  NAND2_X2 U15329 ( .A1(n13347), .A2(n13346), .ZN(n4789) );
  INV_X4 U15330 ( .A(n13414), .ZN(n13349) );
  NAND2_X2 U15331 ( .A1(n13349), .A2(n13348), .ZN(n13355) );
  INV_X4 U15332 ( .A(n13358), .ZN(n13352) );
  INV_X4 U15333 ( .A(n2082), .ZN(n13350) );
  NAND3_X4 U15334 ( .A1(n13352), .A2(n13351), .A3(n13350), .ZN(n13354) );
  NAND2_X2 U15335 ( .A1(n5492), .A2(idOut_20_), .ZN(n13353) );
  OAI211_X2 U15336 ( .C1(ifInst[27]), .C2(n13358), .A(n13357), .B(n13356), 
        .ZN(n13359) );
  INV_X4 U15337 ( .A(n13359), .ZN(n13364) );
  INV_X4 U15338 ( .A(n13360), .ZN(n13362) );
  NAND2_X2 U15339 ( .A1(idOut_29_), .A2(n6589), .ZN(n13361) );
  OAI211_X2 U15340 ( .C1(n13364), .C2(n13363), .A(n13362), .B(n13361), .ZN(
        n4791) );
  INV_X4 U15341 ( .A(n13425), .ZN(n13365) );
  NAND2_X2 U15342 ( .A1(n13365), .A2(n13426), .ZN(n13371) );
  INV_X4 U15343 ( .A(n13366), .ZN(n13368) );
  NAND3_X4 U15344 ( .A1(n13368), .A2(n6581), .A3(n13367), .ZN(n13370) );
  NAND2_X2 U15345 ( .A1(n5492), .A2(idOut_23_), .ZN(n13369) );
  INV_X4 U15346 ( .A(n13372), .ZN(n13376) );
  NAND2_X2 U15347 ( .A1(n5306), .A2(daddr[31]), .ZN(n13374) );
  NAND2_X2 U15348 ( .A1(dwData[31]), .A2(n6609), .ZN(n13373) );
  OAI211_X2 U15349 ( .C1(n13376), .C2(n13375), .A(n13374), .B(n13373), .ZN(
        n13657) );
  NAND2_X2 U15350 ( .A1(ifInst[8]), .A2(n6582), .ZN(n13378) );
  NAND2_X2 U15351 ( .A1(n6587), .A2(aluBoi_imm32w_8_), .ZN(n13377) );
  NAND2_X2 U15352 ( .A1(n13378), .A2(n13377), .ZN(n4802) );
  NAND2_X2 U15353 ( .A1(ifInst[24]), .A2(n6582), .ZN(n13380) );
  NAND2_X2 U15354 ( .A1(n13380), .A2(n13379), .ZN(n13621) );
  NAND2_X2 U15355 ( .A1(ifInst[22]), .A2(n6582), .ZN(n13382) );
  NAND2_X2 U15356 ( .A1(n6587), .A2(net366987), .ZN(n13381) );
  NAND2_X2 U15357 ( .A1(n13382), .A2(n13381), .ZN(n13619) );
  NAND2_X2 U15358 ( .A1(ifInst[20]), .A2(n6582), .ZN(n13384) );
  NAND2_X2 U15359 ( .A1(n6587), .A2(n6835), .ZN(n13383) );
  NAND2_X2 U15360 ( .A1(n13384), .A2(n13383), .ZN(n13617) );
  NAND2_X2 U15361 ( .A1(ifInst[19]), .A2(n6582), .ZN(n13386) );
  NAND2_X2 U15362 ( .A1(n6587), .A2(n6832), .ZN(n13385) );
  NAND2_X2 U15363 ( .A1(n13386), .A2(n13385), .ZN(n13616) );
  NAND2_X2 U15364 ( .A1(ifInst[17]), .A2(n6582), .ZN(n13388) );
  NAND2_X2 U15365 ( .A1(n6804), .A2(n6589), .ZN(n13387) );
  NAND2_X2 U15366 ( .A1(n13388), .A2(n13387), .ZN(n13614) );
  NAND2_X2 U15367 ( .A1(ifInst[15]), .A2(n6582), .ZN(n13420) );
  NAND2_X2 U15368 ( .A1(n6587), .A2(idOut_75_), .ZN(n13389) );
  NAND2_X2 U15369 ( .A1(n13420), .A2(n13389), .ZN(n4808) );
  NAND2_X2 U15370 ( .A1(ifInst[13]), .A2(n6582), .ZN(n13418) );
  NAND2_X2 U15371 ( .A1(n6587), .A2(idOut_73_), .ZN(n13390) );
  NAND2_X2 U15372 ( .A1(n13418), .A2(n13390), .ZN(n4809) );
  NAND2_X2 U15373 ( .A1(ifInst[11]), .A2(n6582), .ZN(n13416) );
  NAND2_X2 U15374 ( .A1(n6587), .A2(idOut_71_), .ZN(n13391) );
  NAND2_X2 U15375 ( .A1(n13416), .A2(n13391), .ZN(n4810) );
  NAND2_X2 U15376 ( .A1(ifInst[6]), .A2(n6582), .ZN(n13393) );
  NAND2_X2 U15377 ( .A1(n6587), .A2(aluBoi_imm32w_6_), .ZN(n13392) );
  NAND2_X2 U15378 ( .A1(n13393), .A2(n13392), .ZN(n13612) );
  NAND2_X2 U15379 ( .A1(ifInst[4]), .A2(n6581), .ZN(n13395) );
  NAND2_X2 U15380 ( .A1(n6587), .A2(aluBoi_imm32w_4_), .ZN(n13394) );
  NAND2_X2 U15381 ( .A1(n13395), .A2(n13394), .ZN(n4812) );
  NAND2_X2 U15382 ( .A1(n6587), .A2(idOut_33_), .ZN(n13397) );
  NAND2_X2 U15383 ( .A1(n13398), .A2(n13397), .ZN(n4813) );
  INV_X4 U15384 ( .A(n13399), .ZN(n13403) );
  MUX2_X2 U15385 ( .A(n13401), .B(n5676), .S(n6586), .Z(n13402) );
  NAND2_X2 U15386 ( .A1(n6587), .A2(n6074), .ZN(n13404) );
  NAND2_X2 U15387 ( .A1(n13405), .A2(n13404), .ZN(n4815) );
  NAND2_X2 U15388 ( .A1(idOut_26_), .A2(n6589), .ZN(n13406) );
  NAND2_X2 U15389 ( .A1(n6587), .A2(aluBoi_imm32w_1_), .ZN(n13407) );
  NAND2_X2 U15390 ( .A1(n13408), .A2(n13407), .ZN(n4817) );
  NAND2_X2 U15391 ( .A1(ifInst[14]), .A2(n6582), .ZN(n13444) );
  NAND2_X2 U15392 ( .A1(n6590), .A2(aluBoi_imm32w_14_), .ZN(n13409) );
  NAND2_X2 U15393 ( .A1(n13444), .A2(n13409), .ZN(n4818) );
  NAND2_X2 U15394 ( .A1(ifInst[12]), .A2(n6581), .ZN(n13442) );
  NAND2_X2 U15395 ( .A1(n6590), .A2(aluBoi_imm32w_12_), .ZN(n13410) );
  NAND2_X2 U15396 ( .A1(n13442), .A2(n13410), .ZN(n4819) );
  NAND2_X2 U15397 ( .A1(ifInst[10]), .A2(n6581), .ZN(n13412) );
  NAND2_X2 U15398 ( .A1(n6590), .A2(aluBoi_imm32w_10_), .ZN(n13411) );
  NAND2_X2 U15399 ( .A1(n13412), .A2(n13411), .ZN(n4820) );
  NAND2_X2 U15400 ( .A1(n13414), .A2(n13413), .ZN(n4821) );
  NAND2_X2 U15401 ( .A1(n6590), .A2(aluBoi_imm32w_11_), .ZN(n13415) );
  NAND2_X2 U15402 ( .A1(n13416), .A2(n13415), .ZN(n4822) );
  NAND2_X2 U15403 ( .A1(n6590), .A2(aluBoi_imm32w_13_), .ZN(n13417) );
  NAND2_X2 U15404 ( .A1(n13418), .A2(n13417), .ZN(n4823) );
  NAND2_X2 U15405 ( .A1(n6590), .A2(aluBoi_imm32w_15_), .ZN(n13419) );
  NAND2_X2 U15406 ( .A1(n13420), .A2(n13419), .ZN(n4824) );
  INV_X4 U15407 ( .A(n13426), .ZN(n13421) );
  NAND3_X4 U15408 ( .A1(n6581), .A2(n13422), .A3(n13421), .ZN(n13424) );
  NAND2_X2 U15409 ( .A1(n6587), .A2(idOut_17_), .ZN(n13423) );
  NAND2_X2 U15410 ( .A1(n13424), .A2(n13423), .ZN(n4825) );
  OAI22_X2 U15411 ( .A1(n5472), .A2(n13430), .B1(n13426), .B2(n13425), .ZN(
        n4826) );
  OAI22_X2 U15412 ( .A1(n5522), .A2(n13430), .B1(n13429), .B2(n13428), .ZN(
        n4828) );
  NAND2_X2 U15413 ( .A1(n5474), .A2(n6582), .ZN(n13432) );
  NAND2_X2 U15414 ( .A1(idOut_34_), .A2(n6589), .ZN(n13431) );
  NAND2_X2 U15415 ( .A1(n13432), .A2(n13431), .ZN(n4829) );
  NOR2_X4 U15416 ( .A1(n13434), .A2(n13433), .ZN(n13501) );
  INV_X4 U15417 ( .A(n13501), .ZN(n13436) );
  NAND2_X2 U15418 ( .A1(idOut_38_), .A2(n6589), .ZN(n13435) );
  NAND2_X2 U15419 ( .A1(n13436), .A2(n13435), .ZN(n4830) );
  NAND2_X2 U15420 ( .A1(ifInst[3]), .A2(n6581), .ZN(n13438) );
  NAND2_X2 U15421 ( .A1(n6590), .A2(aluBoi_imm32w_3_), .ZN(n13437) );
  NAND2_X2 U15422 ( .A1(n13438), .A2(n13437), .ZN(n4831) );
  NAND2_X2 U15423 ( .A1(ifInst[5]), .A2(n6581), .ZN(n13440) );
  NAND2_X2 U15424 ( .A1(n6590), .A2(aluBoi_imm32w_5_), .ZN(n13439) );
  NAND2_X2 U15425 ( .A1(n13440), .A2(n13439), .ZN(n4832) );
  NAND2_X2 U15426 ( .A1(n6588), .A2(idOut_72_), .ZN(n13441) );
  NAND2_X2 U15427 ( .A1(n13442), .A2(n13441), .ZN(n4833) );
  NAND2_X2 U15428 ( .A1(n6587), .A2(idOut_74_), .ZN(n13443) );
  NAND2_X2 U15429 ( .A1(n13444), .A2(n13443), .ZN(n4834) );
  NAND2_X2 U15430 ( .A1(ifInst[16]), .A2(n6581), .ZN(n13446) );
  NAND2_X2 U15431 ( .A1(net369155), .A2(n6590), .ZN(n13445) );
  NAND2_X2 U15432 ( .A1(n13446), .A2(n13445), .ZN(n13613) );
  NAND2_X2 U15433 ( .A1(ifInst[18]), .A2(n6582), .ZN(n13448) );
  NAND2_X2 U15434 ( .A1(n6588), .A2(n6823), .ZN(n13447) );
  NAND2_X2 U15435 ( .A1(n13448), .A2(n13447), .ZN(n13615) );
  NAND2_X2 U15436 ( .A1(ifInst[7]), .A2(n6581), .ZN(n13450) );
  NAND2_X2 U15437 ( .A1(n6590), .A2(aluBoi_imm32w_7_), .ZN(n13449) );
  NAND2_X2 U15438 ( .A1(n13450), .A2(n13449), .ZN(n4837) );
  NAND2_X2 U15439 ( .A1(ifInst[21]), .A2(n6581), .ZN(n13452) );
  NAND2_X2 U15440 ( .A1(n6590), .A2(net367027), .ZN(n13451) );
  NAND2_X2 U15441 ( .A1(n13452), .A2(n13451), .ZN(n13618) );
  NAND2_X2 U15442 ( .A1(ifInst[23]), .A2(n6581), .ZN(n13454) );
  NAND2_X2 U15443 ( .A1(n6590), .A2(net366937), .ZN(n13453) );
  NAND2_X2 U15444 ( .A1(n13454), .A2(n13453), .ZN(n13620) );
  NAND2_X2 U15445 ( .A1(n5313), .A2(n6581), .ZN(n13456) );
  NAND2_X2 U15446 ( .A1(n6590), .A2(n6787), .ZN(n13455) );
  NAND2_X2 U15447 ( .A1(n13456), .A2(n13455), .ZN(n13622) );
  NAND2_X2 U15448 ( .A1(ifInst[9]), .A2(n6583), .ZN(n13458) );
  NAND2_X2 U15449 ( .A1(n6590), .A2(aluBoi_imm32w_9_), .ZN(n13457) );
  NAND2_X2 U15450 ( .A1(n13458), .A2(n13457), .ZN(n4841) );
  INV_X4 U15451 ( .A(inst[0]), .ZN(n13459) );
  INV_X4 U15452 ( .A(inst[1]), .ZN(n13460) );
  OAI22_X2 U15453 ( .A1(n6602), .A2(n13460), .B1(n6594), .B2(n13499), .ZN(
        n13577) );
  INV_X4 U15454 ( .A(inst[2]), .ZN(n13461) );
  INV_X4 U15455 ( .A(inst[3]), .ZN(n13462) );
  OAI22_X2 U15456 ( .A1(n6602), .A2(n13462), .B1(n6594), .B2(n5343), .ZN(
        n13579) );
  INV_X4 U15457 ( .A(inst[4]), .ZN(n13463) );
  OAI22_X2 U15458 ( .A1(n6602), .A2(n13463), .B1(n6594), .B2(n5456), .ZN(
        n13580) );
  INV_X4 U15459 ( .A(inst[5]), .ZN(n13464) );
  OAI22_X2 U15460 ( .A1(n6602), .A2(n13464), .B1(n6594), .B2(n5346), .ZN(
        n13581) );
  INV_X4 U15461 ( .A(inst[6]), .ZN(n13465) );
  OAI22_X2 U15462 ( .A1(n6602), .A2(n13465), .B1(n6594), .B2(n5464), .ZN(
        n13582) );
  INV_X4 U15463 ( .A(inst[7]), .ZN(n13466) );
  OAI22_X2 U15464 ( .A1(n6602), .A2(n13466), .B1(n6594), .B2(n5480), .ZN(
        n13583) );
  INV_X4 U15465 ( .A(inst[8]), .ZN(n13467) );
  OAI22_X2 U15466 ( .A1(n6602), .A2(n13467), .B1(n6594), .B2(n5469), .ZN(
        n13584) );
  INV_X4 U15467 ( .A(inst[9]), .ZN(n13468) );
  OAI22_X2 U15468 ( .A1(n6602), .A2(n13468), .B1(n6594), .B2(n5481), .ZN(
        n13585) );
  INV_X4 U15469 ( .A(inst[10]), .ZN(n13469) );
  OAI22_X2 U15470 ( .A1(n6602), .A2(n13469), .B1(n6595), .B2(n5465), .ZN(
        n13586) );
  INV_X4 U15471 ( .A(inst[11]), .ZN(n13470) );
  OAI22_X2 U15472 ( .A1(n6602), .A2(n13470), .B1(n6595), .B2(n5475), .ZN(
        n13587) );
  INV_X4 U15473 ( .A(inst[12]), .ZN(n13471) );
  OAI22_X2 U15474 ( .A1(n6602), .A2(n13471), .B1(n6595), .B2(n5463), .ZN(
        n13588) );
  INV_X4 U15475 ( .A(inst[13]), .ZN(n13472) );
  OAI22_X2 U15476 ( .A1(n6602), .A2(n13472), .B1(n6595), .B2(n5473), .ZN(
        n13589) );
  INV_X4 U15477 ( .A(inst[14]), .ZN(n13473) );
  OAI22_X2 U15478 ( .A1(n6602), .A2(n13473), .B1(n6595), .B2(n5468), .ZN(
        n13590) );
  INV_X4 U15479 ( .A(inst[15]), .ZN(n13474) );
  OAI22_X2 U15480 ( .A1(n6602), .A2(n13474), .B1(n6595), .B2(n5485), .ZN(
        n13591) );
  INV_X4 U15481 ( .A(inst[16]), .ZN(n13475) );
  OAI22_X2 U15482 ( .A1(n6602), .A2(n13475), .B1(n6595), .B2(n5467), .ZN(
        n13592) );
  INV_X4 U15483 ( .A(inst[17]), .ZN(n13476) );
  OAI22_X2 U15484 ( .A1(n6601), .A2(n13476), .B1(n6595), .B2(n5493), .ZN(
        n13593) );
  INV_X4 U15485 ( .A(inst[18]), .ZN(n13477) );
  OAI22_X2 U15486 ( .A1(n6601), .A2(n13477), .B1(n6595), .B2(n5479), .ZN(
        n13594) );
  INV_X4 U15487 ( .A(inst[19]), .ZN(n13478) );
  OAI22_X2 U15488 ( .A1(n6601), .A2(n13478), .B1(n6595), .B2(n5494), .ZN(
        n13595) );
  INV_X4 U15489 ( .A(inst[20]), .ZN(n13479) );
  OAI22_X2 U15490 ( .A1(n6601), .A2(n13479), .B1(n6595), .B2(n5470), .ZN(
        n13596) );
  INV_X4 U15491 ( .A(inst[21]), .ZN(n13481) );
  INV_X4 U15492 ( .A(ifInst[21]), .ZN(n13480) );
  OAI22_X2 U15493 ( .A1(n6601), .A2(n13481), .B1(n6594), .B2(n13480), .ZN(
        n13597) );
  INV_X4 U15494 ( .A(inst[22]), .ZN(n13483) );
  INV_X4 U15495 ( .A(ifInst[22]), .ZN(n13482) );
  OAI22_X2 U15496 ( .A1(n6601), .A2(n13483), .B1(n6594), .B2(n13482), .ZN(
        n13598) );
  INV_X4 U15497 ( .A(inst[23]), .ZN(n13485) );
  INV_X4 U15498 ( .A(ifInst[23]), .ZN(n13484) );
  OAI22_X2 U15499 ( .A1(n6601), .A2(n13485), .B1(n6594), .B2(n13484), .ZN(
        n13599) );
  INV_X4 U15500 ( .A(inst[24]), .ZN(n13487) );
  INV_X4 U15501 ( .A(ifInst[24]), .ZN(n13486) );
  OAI22_X2 U15502 ( .A1(n6601), .A2(n13487), .B1(n6594), .B2(n13486), .ZN(
        n13600) );
  INV_X4 U15503 ( .A(inst[25]), .ZN(n13489) );
  OAI22_X2 U15504 ( .A1(n6601), .A2(n13489), .B1(n6594), .B2(n13488), .ZN(
        n13601) );
  INV_X4 U15505 ( .A(inst[26]), .ZN(n13490) );
  OAI22_X2 U15506 ( .A1(n6601), .A2(n13490), .B1(n13539), .B2(n6594), .ZN(
        n13602) );
  INV_X4 U15507 ( .A(inst[27]), .ZN(n13492) );
  OAI22_X2 U15508 ( .A1(n6601), .A2(n13492), .B1(n13491), .B2(n6594), .ZN(
        n13603) );
  INV_X4 U15509 ( .A(inst[28]), .ZN(n13494) );
  OAI22_X2 U15510 ( .A1(n6601), .A2(n13494), .B1(n6594), .B2(n13493), .ZN(
        n13604) );
  INV_X4 U15511 ( .A(inst[29]), .ZN(n13496) );
  OAI22_X2 U15512 ( .A1(n6601), .A2(n13496), .B1(n6594), .B2(n13495), .ZN(
        n13605) );
  INV_X4 U15513 ( .A(inst[31]), .ZN(n13498) );
  OAI22_X2 U15514 ( .A1(n6601), .A2(n13498), .B1(n13497), .B2(n6594), .ZN(
        n13607) );
  XOR2_X2 U15515 ( .A(ifInst[3]), .B(ifInst[4]), .Z(n13502) );
  NAND4_X2 U15516 ( .A1(n13503), .A2(n13502), .A3(n13501), .A4(n13500), .ZN(
        n13505) );
  NAND2_X2 U15517 ( .A1(n6588), .A2(didMult), .ZN(n13504) );
  NAND2_X2 U15518 ( .A1(n13505), .A2(n13504), .ZN(n4874) );
  INV_X4 U15519 ( .A(inst[30]), .ZN(n13507) );
  OAI22_X2 U15520 ( .A1(n6602), .A2(n13507), .B1(n6594), .B2(n5455), .ZN(
        n13606) );
  NAND2_X2 U15521 ( .A1(n6609), .A2(daddr[31]), .ZN(n13518) );
  AOI22_X2 U15522 ( .A1(aluBoi_multBoi_temppp[28]), .A2(net368069), .B1(n5316), 
        .B2(aluBoi_imm32w_15_), .ZN(n13517) );
  OAI21_X4 U15523 ( .B1(n13513), .B2(n13512), .A(n13062), .ZN(n13516) );
  NAND4_X2 U15524 ( .A1(n13515), .A2(n13517), .A3(n13516), .A4(n13518), .ZN(
        n4876) );
  INV_X4 U15525 ( .A(n3391), .ZN(n13662) );
  INV_X4 U15526 ( .A(n3083), .ZN(n13663) );
  INV_X4 U15527 ( .A(n2992), .ZN(n13664) );
  INV_X4 U15528 ( .A(n2991), .ZN(n13665) );
  INV_X4 U15529 ( .A(n2990), .ZN(n13666) );
  INV_X4 U15530 ( .A(n2989), .ZN(n13667) );
  INV_X4 U15531 ( .A(n2988), .ZN(n13668) );
  INV_X4 U15532 ( .A(n2987), .ZN(n13669) );
  INV_X4 U15533 ( .A(n2986), .ZN(n13670) );
  INV_X4 U15534 ( .A(n2984), .ZN(n13671) );
  INV_X4 U15535 ( .A(n2983), .ZN(n13672) );
  INV_X4 U15536 ( .A(n1213), .ZN(n13674) );
  INV_X4 U15537 ( .A(drData[15]), .ZN(n13676) );
  INV_X4 U15538 ( .A(n1232), .ZN(n13677) );
  NOR2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U218 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n14), .A2(n6606), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n107) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U217 ( .A1(n6545), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(net377611), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n185) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U216 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n49), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n44), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n185), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n184) );
  NAND2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U215 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n102) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U214 ( .A1(n5231), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .B2(n6521), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n183) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U213 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n32), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n65), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n183), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n86) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U212 ( .A1(n6527), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6529), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n182) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U211 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n35), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n63), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n182), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n85) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U210 ( .A1(n6511), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6513), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n181) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U209 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n70), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n20), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n181), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n126) );
  AND2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U208 ( .A1(n6616), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n15), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n133) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U207 ( .A1(n6517), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n5309), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n180) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U206 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n29), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n68), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n180), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n127) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U205 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n148), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n126), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n127), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n179) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U204 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n86), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n85), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n18), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n150) );
  AND2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U203 ( .A1(n6616), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n16), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n176) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U202 ( .A1(n6535), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6537), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n178) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U201 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n60), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n61), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n178), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n84) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U200 ( .A1(net368498), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(net345751), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n177) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U199 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n47), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n46), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n177), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n174) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U198 ( .A1(n13706), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n10770), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n175) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U197 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n52), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n55), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n175), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n87) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U196 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n84), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n71), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n174), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n87), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n173) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U195 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n43), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n102), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n150), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n173), .ZN(aluBoi_aluBoi_shft_sraout[0])
         );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U194 ( .A1(n6539), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(net368519), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n172) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U193 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n56), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n59), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n172), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n95) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U192 ( .A1(n6515), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(net368584), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n171) );
  NAND2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U191 ( .A1(
        aluBoi_aluBoi_shft_sraout[31]), .A2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n146) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U190 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n134), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n130), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n23), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n122) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U189 ( .A1(n13527), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6533), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n170) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U188 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n62), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n37), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n170), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n96) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U187 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .A2(n6523), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .B2(n6525), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n169) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U186 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n64), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n33), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n169), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n97) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U185 ( .A1(net377607), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(net368572), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n168) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U184 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n66), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n30), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n168), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n131) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U183 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n96), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n97), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n131), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n167) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U182 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n51), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n122), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n167), .ZN(aluBoi_aluBoi_shft_sraout[10]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U181 ( .A1(n6537), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6539), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n166) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U180 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n59), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n60), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n166), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n90) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U179 ( .A1(n6513), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6515), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n165) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U178 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n69), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n70), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n165), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n128) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U177 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n15), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n20), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n146), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n153) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U176 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n128), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n153), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n121) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U175 ( .A1(n6529), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n13527), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n164) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U174 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n37), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n35), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n164), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n91) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U173 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .A2(n6521), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .B2(n6523), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n163) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U172 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n33), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n32), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n163), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n92) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U171 ( .A1(n5309), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(net377607), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n162) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U170 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n30), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n29), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n162), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n129) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U169 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n91), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n92), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n129), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n161) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U168 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n54), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n121), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n161), .ZN(aluBoi_aluBoi_shft_sraout[11]) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U167 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n126), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n153), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n120) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U166 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n85), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n86), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n127), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n160) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U165 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n57), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n120), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n160), .ZN(aluBoi_aluBoi_shft_sraout[12]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U164 ( .A1(n6533), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n6535), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n159) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U163 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n61), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n62), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n159), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n76) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U162 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .A2(n6511), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B2(n6509), .C1(n6606), .C2(
        aluBoi_aluBoi_shft_sraout[31]), .ZN(aluBoi_aluBoi_shft_SRA_sra_25_n158) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U161 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n27), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n153), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n119) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U160 ( .A1(n6525), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(n6527), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n157) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U159 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n63), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n64), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n157), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n78) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U158 ( .A1(net368572), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n5231), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n156) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U157 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n65), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n66), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n156), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n80) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U156 ( .A1(net368584), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(n6517), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n108), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n155) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U155 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n6), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n68), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n67), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n155), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n124) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U154 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n78), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n80), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n124), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n154) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U153 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n58), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n119), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n154), .ZN(aluBoi_aluBoi_shft_sraout[13]) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U152 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n134), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n153), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n111) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U151 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n97), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n131), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n130), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n152) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U150 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n36), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n111), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n152), .ZN(aluBoi_aluBoi_shft_sraout[14]) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U149 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n128), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n129), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n28), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n151) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U148 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n31), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n102), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n34), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n151), .ZN(aluBoi_aluBoi_shft_sraout[15]) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U147 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n150), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[16]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U146 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n148), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n27), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n124), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n149) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U145 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n80), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n78), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n26), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n138) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U144 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n138), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[17]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U143 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n148), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n134), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n130), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n147) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U142 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n131), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n97), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n21), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n113) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U141 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n113), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[18]) );
  NOR2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U140 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n146), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n15), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n135) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U139 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n128), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n135), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n145) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U138 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n129), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n92), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n24), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n103) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U137 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n103), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[19]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U136 ( .A1(n6543), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(n6545), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n144) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U135 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n44), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n41), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n144), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n143) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U134 ( .A1(net368502), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(net368498), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n142) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U133 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n46), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n45), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n142), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n140) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U132 ( .A1(net368519), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(n13706), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n141) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U131 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n55), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n56), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n141), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n81) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U130 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n76), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n71), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n140), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n81), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n139) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U129 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n39), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n102), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n138), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n139), .ZN(aluBoi_aluBoi_shft_sraout[1])
         );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U128 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n126), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n135), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n137) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U127 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n127), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n86), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n19), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n100) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U126 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n100), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[20]) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U125 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n27), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n135), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n136) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U124 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n124), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n80), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n25), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n98) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U123 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n98), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[21]) );
  AOI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U122 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n133), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n134), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n135), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n132) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U121 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n93), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[22]) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U120 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n128), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n129), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n23), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n88) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U119 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n88), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[23]) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U118 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n126), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n127), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n23), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n82) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U117 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n82), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[24]) );
  AOI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U116 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n27), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n124), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n23), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n74) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U115 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n74), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[25]) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U114 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n122), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[26]) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U113 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n121), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[27]) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U112 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n120), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[28]) );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U111 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n119), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[29]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U110 ( .A1(n6541), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(n6543), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n118) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U109 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n41), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n53), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n118), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n117) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U108 ( .A1(n13525), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(net368502), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n116) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U107 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n45), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n48), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n116), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n115) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U106 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n96), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n71), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n115), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n95), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n114) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U105 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n40), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n102), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n113), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n114), .ZN(aluBoi_aluBoi_shft_sraout[2])
         );
  OAI21_X1 aluBoi_aluBoi_shft_SRA_sra_25_U104 ( .B1(n6618), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n111), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(aluBoi_aluBoi_shft_sraout[30]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U103 ( .A1(n10770), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n9), .B1(n6541), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n110) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U102 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n53), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n7), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n52), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n110), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n109) );
  AOI22_X1 aluBoi_aluBoi_shft_SRA_sra_25_U101 ( .A1(net377611), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n10), .B1(n13525), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n12), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n106) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U100 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n48), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n49), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n106), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n105) );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U99 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n91), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n71), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n105), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n90), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n104) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U98 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n38), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n102), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n103), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n104), .ZN(aluBoi_aluBoi_shft_sraout[3])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U97 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n87), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n84), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n85), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n101) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U96 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n43), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n100), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n101), .ZN(aluBoi_aluBoi_shft_sraout[4])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U95 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n81), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n76), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n78), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n99) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U94 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n39), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n98), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n99), .ZN(aluBoi_aluBoi_shft_sraout[5])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U93 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n95), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n96), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n97), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n94) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U92 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n40), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n93), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n94), .ZN(aluBoi_aluBoi_shft_sraout[6])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U91 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n90), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n91), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n92), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n89) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U90 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n38), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n88), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n89), .ZN(aluBoi_aluBoi_shft_sraout[7])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U89 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n84), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n85), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n86), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n83) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U88 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n42), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n82), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n83), .ZN(aluBoi_aluBoi_shft_sraout[8])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRA_sra_25_U87 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n72), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n76), .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n77), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n78), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n79), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n80), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n75) );
  OAI221_X1 aluBoi_aluBoi_shft_SRA_sra_25_U86 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n50), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n74), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n75), .ZN(aluBoi_aluBoi_shft_sraout[9])
         );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U85 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n73), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n71) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U84 ( .A(n6509), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n70) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U83 ( .A(n6515), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n68) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U82 ( .A(n6513), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n67) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U81 ( .A(n5309), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n66) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U80 ( .A(n6521), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n64) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U79 ( .A(n6523), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n63) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U78 ( .A(n6529), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n62) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U77 ( .A(n13527), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n61) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U76 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n76), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n58) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U75 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n84), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n57) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U74 ( .A(n6537), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n56) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U73 ( .A(n6539), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n55) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U72 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n90), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n54) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U71 ( .A(n13706), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n53) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U70 ( .A(net368519), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n52) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U69 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n95), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n51) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U68 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n81), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n50) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U67 ( .A(n6543), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n49) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U66 ( .A(n6545), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n48) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U65 ( .A(net368502), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n47) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U64 ( .A(n13525), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n46) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U63 ( .A(n6541), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n44) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U62 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n184), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n43) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U61 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n87), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n42) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U60 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n117), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n40) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U59 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n143), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n39) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U58 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n109), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n38) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U57 ( .A(n6527), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n37) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U56 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n96), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n36) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U55 ( .A(n6525), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n35) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U54 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n91), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n34) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U53 ( .A(net368572), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n32) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U52 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n92), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n31) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U51 ( .A(n6517), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n30) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U50 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n112), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n28) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U49 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n158), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n27) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U48 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n149), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n26) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U47 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n136), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n25) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U46 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n145), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n24) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U45 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n146), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n23) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U44 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n147), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n21) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U43 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n137), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n19) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U42 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n179), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n18) );
  INV_X32 aluBoi_aluBoi_shft_SRA_sra_25_U41 ( .A(n6618), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n17) );
  NOR2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U40 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n15), .A2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n123) );
  NOR2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U39 ( .A1(n6614), .A2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n125) );
  INV_X32 aluBoi_aluBoi_shft_SRA_sra_25_U38 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n3), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n4) );
  AND2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U37 ( .A1(n6614), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n176), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n79) );
  NAND2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U36 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n17), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n73) );
  AND2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U35 ( .A1(
        aluBoi_aluBoi_shft_SRA_sra_25_n176), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n15), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n77) );
  INV_X8 aluBoi_aluBoi_shft_SRA_sra_25_U34 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n102), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n72) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U33 ( .A(n10770), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n41) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U32 ( .A(n6511), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n69) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U31 ( .A(net377607), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n65) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U30 ( .A(n5231), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n33) );
  INV_X1 aluBoi_aluBoi_shft_SRA_sra_25_U29 ( .A(n6535), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n59) );
  INV_X1 aluBoi_aluBoi_shft_SRA_sra_25_U28 ( .A(n6533), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n60) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U27 ( .A(net377611), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n45) );
  INV_X1 aluBoi_aluBoi_shft_SRA_sra_25_U26 ( .A(net368584), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n29) );
  AND2_X2 aluBoi_aluBoi_shft_SRA_sra_25_U25 ( .A1(n6614), .A2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n148) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U24 ( .A(n6614), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n15) );
  OAI221_X2 aluBoi_aluBoi_shft_SRA_sra_25_U23 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n5), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n67), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n8), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n69), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n171), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n130) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U22 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n132), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n22) );
  AOI221_X2 aluBoi_aluBoi_shft_SRA_sra_25_U21 ( .B1(
        aluBoi_aluBoi_shft_SRA_sra_25_n130), .B2(
        aluBoi_aluBoi_shft_SRA_sra_25_n123), .C1(
        aluBoi_aluBoi_shft_SRA_sra_25_n131), .C2(
        aluBoi_aluBoi_shft_SRA_sra_25_n4), .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n22), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n93) );
  NOR2_X2 aluBoi_aluBoi_shft_SRA_sra_25_U20 ( .A1(n6612), .A2(n6606), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n108) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U19 ( .A(n6612), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n14) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U18 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n2), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n5) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U17 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n11), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n10) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U16 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n107), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n11) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U15 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n1), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n8) );
  INV_X8 aluBoi_aluBoi_shft_SRA_sra_25_U14 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n13), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n12) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U13 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n108), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n13) );
  AND2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U12 ( .A1(n6606), .A2(
        aluBoi_aluBoi_shft_SRA_sra_25_n14), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n2) );
  AND2_X4 aluBoi_aluBoi_shft_SRA_sra_25_U11 ( .A1(n6612), .A2(n6606), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n1) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U10 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n125), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n3) );
  INV_X8 aluBoi_aluBoi_shft_SRA_sra_25_U9 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n1), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n7) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U8 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n11), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n9) );
  INV_X4 aluBoi_aluBoi_shft_SRA_sra_25_U7 ( .A(
        aluBoi_aluBoi_shft_SRA_sra_25_n2), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n6) );
  MUX2_X2 aluBoi_aluBoi_shft_SRA_sra_25_U6 ( .A(aluBoi_aluBoi_shft_sraout[31]), 
        .B(n6509), .S(aluBoi_aluBoi_shft_SRA_sra_25_n108), .Z(
        aluBoi_aluBoi_shft_SRA_sra_25_n134) );
  INV_X2 aluBoi_aluBoi_shft_SRA_sra_25_U5 ( .A(aluBoi_aluBoi_shft_sraout[31]), 
        .ZN(aluBoi_aluBoi_shft_SRA_sra_25_n20) );
  NAND2_X1 aluBoi_aluBoi_shft_SRA_sra_25_U4 ( .A1(n6618), .A2(
        aluBoi_aluBoi_shft_sraout[31]), .ZN(aluBoi_aluBoi_shft_SRA_sra_25_n112) );
  INV_X1 aluBoi_aluBoi_shft_SRA_sra_25_U3 ( .A(n6618), .ZN(
        aluBoi_aluBoi_shft_SRA_sra_25_n16) );
  NAND2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U215 ( .A1(n6606), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n16), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n109) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U214 ( .A1(n6545), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(net377611), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n184) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U213 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n47), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n52), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n184), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n183) );
  NAND2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U212 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n103) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U211 ( .A1(n6519), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .B2(n6521), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n182) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U210 ( .A1(n6527), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(n6529), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n181) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U209 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n64), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n39), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n181), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n86) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U208 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n17), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n18), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n144) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U207 ( .A1(n6511), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(n6513), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n180) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U206 ( .A1(n6517), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(n5309), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n179) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U205 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n69), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n33), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n179), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n129) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U204 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n144), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n124), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n129), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n178) );
  AOI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U203 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n87), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n86), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n22), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n146) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U202 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n18), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n19), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n175) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U201 ( .A1(n6535), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(n6537), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n177) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U200 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n62), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n61), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n177), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n85) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U199 ( .A1(net368498), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(net345751), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n176) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U198 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n49), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n50), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n176), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n173) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U197 ( .A1(n13706), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n8), .B1(n10724), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n174) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U196 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n58), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n55), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n174), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n88) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U195 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n85), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n173), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n88), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n172) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U194 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n46), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n146), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n172), .ZN(aluBoi_aluBoi_shft_srlout[0])
         );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U193 ( .A1(n6539), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(net368519), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n171) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U192 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n60), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n59), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n171), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n96) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U191 ( .A1(n6515), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(net368584), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n170) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U190 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n70), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n68), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n170), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n133) );
  OAI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U189 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n12), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n71), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n9), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n32), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n116) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U188 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n133), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n116), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n125) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U187 ( .A1(n13527), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6533), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n169) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U186 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n40), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n63), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n169), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n97) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U185 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .A2(n6523), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .B2(n6525), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n168) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U184 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n37), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n65), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n168), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n98) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U183 ( .A1(net377607), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n111), .B1(net368572), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n167) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U182 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n97), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n98), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n134), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n166) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U181 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n54), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n125), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n166), .ZN(aluBoi_aluBoi_shft_srlout[10]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U180 ( .A1(n6529), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n13527), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n165) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U179 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n39), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n40), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n165), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n92) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U178 ( .A1(n6537), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6539), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n164) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U177 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n61), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n60), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n164), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n91) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U176 ( .A1(n5309), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(net377607), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n163) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U175 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n33), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n34), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n163), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n132) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U174 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n32), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n12), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n115) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U173 ( .A1(n6513), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n111), .B1(n6515), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n162) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U172 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .A2(n6521), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .B2(n6523), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n161) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U171 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n36), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n37), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n161), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n93) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U170 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n132), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n160), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n93), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n159) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U169 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n38), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n57), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n159), .ZN(aluBoi_aluBoi_shft_srlout[11]) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U168 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n129), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n148), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n124), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n87), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n158) );
  AOI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U167 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n86), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n85), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n24), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n157) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U166 ( .A1(n6525), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6527), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n156) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U165 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n65), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n64), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n156), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n79) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U164 ( .A1(n6533), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6535), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n155) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U163 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n63), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n62), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n155), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n77) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U162 ( .A1(net368584), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6517), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n154) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U161 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n68), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n69), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n154), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n126) );
  OAI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U160 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n9), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n71), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n32), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n12), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n70), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n123) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U159 ( .A1(net368572), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6519), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n153) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U158 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n67), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n66), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n153), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n81) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U157 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n126), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n148), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n123), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n81), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n152) );
  AOI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U156 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n79), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n77), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n30), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n151) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U155 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n133), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n148), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n116), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n134), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n150) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U154 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n130), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n148), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n115), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n132), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n147) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U153 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n35), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n38), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n147), .ZN(aluBoi_aluBoi_shft_srlout[15]) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U152 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n146), .ZN(aluBoi_aluBoi_shft_srlout[16]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U151 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n144), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n123), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n126), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n145) );
  AOI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U150 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n81), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n79), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n31), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n135) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U149 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n135), .ZN(aluBoi_aluBoi_shft_srlout[17]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U148 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n144), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n116), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n133), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n143) );
  AOI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U147 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n134), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n98), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n27), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n117) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U146 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n117), .ZN(aluBoi_aluBoi_shft_srlout[18]) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U145 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n93), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n132), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n142), .C2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n104) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U144 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n104), .ZN(aluBoi_aluBoi_shft_srlout[19]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U143 ( .A1(n6543), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6545), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n141) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U142 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n44), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n47), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n141), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n140) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U141 ( .A1(net376602), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(net368498), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n139) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U140 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n48), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n49), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n139), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n137) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U139 ( .A1(net368519), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n13706), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n138) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U138 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n59), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n58), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n138), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n82) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U137 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n77), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n137), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n82), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n136) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U136 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n42), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n135), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n136), .ZN(aluBoi_aluBoi_shft_srlout[1])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U135 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n129), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n124), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n87), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n101) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U134 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n101), .ZN(aluBoi_aluBoi_shft_srlout[20]) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U133 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n126), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n123), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n81), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n99) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U132 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n99), .ZN(aluBoi_aluBoi_shft_srlout[21])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U131 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n133), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n116), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n134), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n94) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U130 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n94), .ZN(aluBoi_aluBoi_shft_srlout[22])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U129 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n130), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n115), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n131), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n132), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n89) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U128 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n89), .ZN(aluBoi_aluBoi_shft_srlout[23])
         );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U127 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n129), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n124), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n83) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U126 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n83), .ZN(aluBoi_aluBoi_shft_srlout[24])
         );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U125 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n126), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n123), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n128), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n75) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U124 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n75), .ZN(aluBoi_aluBoi_shft_srlout[25])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U123 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n125), .ZN(aluBoi_aluBoi_shft_srlout[26]) );
  NOR3_X1 aluBoi_aluBoi_shft_SRL_srl_16_U122 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n28), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .A3(n6616), .ZN(
        aluBoi_aluBoi_shft_srlout[27]) );
  AND2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U121 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n124), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .ZN(aluBoi_aluBoi_shft_srlout[28]) );
  AND2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U120 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n123), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .ZN(aluBoi_aluBoi_shft_srlout[29]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U119 ( .A1(n6541), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6543), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n122) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U118 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n56), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n44), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n122), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n121) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U117 ( .A1(n13525), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(net376602), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n120) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U116 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n51), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n48), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n120), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n119) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U115 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n97), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n119), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n96), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n118) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U114 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n43), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n117), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n118), .ZN(aluBoi_aluBoi_shft_srlout[2])
         );
  AND2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U113 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n116), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .ZN(aluBoi_aluBoi_shft_srlout[30]) );
  AND2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U112 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n115), .ZN(aluBoi_aluBoi_shft_srlout[31]) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U111 ( .A1(n10724), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n6541), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n13), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n114) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U110 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n55), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n56), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n114), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n113) );
  AOI22_X1 aluBoi_aluBoi_shft_SRL_srl_16_U109 ( .A1(net377611), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n7), .B1(n13525), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n14), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n110) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U108 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n52), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n51), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n110), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n107) );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U107 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n92), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n107), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n91), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n105) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U106 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n41), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n104), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n105), .ZN(aluBoi_aluBoi_shft_srlout[3])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U105 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n88), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n85), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n86), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n102) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U104 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n46), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n101), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n102), .ZN(aluBoi_aluBoi_shft_srlout[4])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U103 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n82), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n77), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n79), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n100) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U102 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n42), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n99), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n100), .ZN(aluBoi_aluBoi_shft_srlout[5])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U101 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n96), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n97), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n98), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n95) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U100 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n43), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n94), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n95), .ZN(aluBoi_aluBoi_shft_srlout[6])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U99 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n91), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n92), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n93), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n90) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U98 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n41), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n89), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n90), .ZN(aluBoi_aluBoi_shft_srlout[7])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U97 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n85), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n86), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n87), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n84) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U96 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n45), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n83), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n84), .ZN(aluBoi_aluBoi_shft_srlout[8])
         );
  AOI222_X1 aluBoi_aluBoi_shft_SRL_srl_16_U95 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n77), .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n78), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n79), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n80), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n81), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n76) );
  OAI221_X1 aluBoi_aluBoi_shft_SRL_srl_16_U94 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n53), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n72), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n75), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n76), .ZN(aluBoi_aluBoi_shft_srlout[9])
         );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U93 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n127), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n73) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U92 ( .A(n6509), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n71) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U91 ( .A(n6515), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n69) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U90 ( .A(n6513), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n68) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U89 ( .A(n5309), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n67) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U88 ( .A(n6521), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n65) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U87 ( .A(n6523), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n64) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U86 ( .A(n6529), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n63) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U85 ( .A(n13527), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n62) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U84 ( .A(n6537), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n59) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U83 ( .A(n6539), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n58) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U82 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n91), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n57) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U81 ( .A(n13706), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n56) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U80 ( .A(net368519), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n55) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U79 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n96), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n54) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U78 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n82), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n53) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U77 ( .A(n6543), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n52) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U76 ( .A(n6545), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n51) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U75 ( .A(net376602), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n50) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U74 ( .A(n13525), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n49) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U73 ( .A(net377611), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n48) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U72 ( .A(n6541), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n47) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U71 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n183), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n46) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U70 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n88), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n45) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U69 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n121), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n43) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U68 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n140), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n42) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U67 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n113), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n41) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U66 ( .A(n6527), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n40) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U65 ( .A(n6525), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n39) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U64 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n92), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n38) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U63 ( .A(net368572), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n36) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U62 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n93), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n35) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U61 ( .A(n6517), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n34) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U60 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n145), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n31) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U59 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n152), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n30) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U58 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n151), .ZN(aluBoi_aluBoi_shft_srlout[13]) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U57 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n142), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n28) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U56 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n143), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n27) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U55 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n149), .ZN(aluBoi_aluBoi_shft_srlout[14]) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U54 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n158), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n24) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U53 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n157), .ZN(aluBoi_aluBoi_shft_srlout[12]) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U52 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n178), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n22) );
  INV_X32 aluBoi_aluBoi_shft_SRL_srl_16_U51 ( .A(n6618), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n20) );
  INV_X16 aluBoi_aluBoi_shft_SRL_srl_16_U50 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n11), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n15) );
  INV_X32 aluBoi_aluBoi_shft_SRL_srl_16_U49 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n15), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n14) );
  INV_X32 aluBoi_aluBoi_shft_SRL_srl_16_U48 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n15), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n13) );
  INV_X16 aluBoi_aluBoi_shft_SRL_srl_16_U47 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n111), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n10) );
  INV_X32 aluBoi_aluBoi_shft_SRL_srl_16_U46 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n3), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n1) );
  NOR2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U45 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n17), .A2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n128) );
  AND2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U44 ( .A1(n6614), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n175), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n80) );
  NOR2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U43 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n73), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n21), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n106) );
  AND2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U42 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n175), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n17), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n78) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U41 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n103), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n74) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U40 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n72) );
  INV_X2 aluBoi_aluBoi_shft_SRL_srl_16_U39 ( .A(n10724), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n44) );
  INV_X2 aluBoi_aluBoi_shft_SRL_srl_16_U38 ( .A(n6511), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n70) );
  INV_X2 aluBoi_aluBoi_shft_SRL_srl_16_U37 ( .A(net377607), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n66) );
  INV_X2 aluBoi_aluBoi_shft_SRL_srl_16_U36 ( .A(n6519), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n37) );
  INV_X1 aluBoi_aluBoi_shft_SRL_srl_16_U35 ( .A(n6535), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n60) );
  INV_X1 aluBoi_aluBoi_shft_SRL_srl_16_U34 ( .A(n6533), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n61) );
  INV_X1 aluBoi_aluBoi_shft_SRL_srl_16_U33 ( .A(net368584), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n33) );
  NOR2_X2 aluBoi_aluBoi_shft_SRL_srl_16_U32 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n18), .A2(n6614), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n131) );
  NOR2_X1 aluBoi_aluBoi_shft_SRL_srl_16_U31 ( .A1(n6614), .A2(n6616), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n127) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U30 ( .A(n6614), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n17) );
  OAI221_X2 aluBoi_aluBoi_shft_SRL_srl_16_U29 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n34), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n67), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n167), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n134) );
  NOR2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U28 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n16), .A2(n6606), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n111) );
  OAI221_X2 aluBoi_aluBoi_shft_SRL_srl_16_U27 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n2), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n71), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n5), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n70), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n162), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n130) );
  MUX2_X2 aluBoi_aluBoi_shft_SRL_srl_16_U26 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n115), .B(
        aluBoi_aluBoi_shft_SRL_srl_16_n130), .S(
        aluBoi_aluBoi_shft_SRL_srl_16_n17), .Z(
        aluBoi_aluBoi_shft_SRL_srl_16_n142) );
  NOR2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U25 ( .A1(n6612), .A2(n6606), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n112) );
  NAND2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U24 ( .A1(n6606), .A2(n6612), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n108) );
  INV_X2 aluBoi_aluBoi_shft_SRL_srl_16_U23 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n150), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n26) );
  AOI221_X2 aluBoi_aluBoi_shft_SRL_srl_16_U22 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n98), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n74), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n97), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n106), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n26), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n149) );
  NOR2_X4 aluBoi_aluBoi_shft_SRL_srl_16_U21 ( .A1(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n73), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n148) );
  OAI221_X2 aluBoi_aluBoi_shft_SRL_srl_16_U20 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n66), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n36), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n182), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n87) );
  NOR2_X2 aluBoi_aluBoi_shft_SRL_srl_16_U19 ( .A1(n6616), .A2(
        aluBoi_aluBoi_shft_SRL_srl_16_n28), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n160) );
  INV_X16 aluBoi_aluBoi_shft_SRL_srl_16_U18 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n10), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n7) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U17 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n6), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n4) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U16 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n109), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n6) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U15 ( .A(n6616), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n18) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U14 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n112), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n12) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U13 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n12), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n11) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U12 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n19) );
  OAI221_X2 aluBoi_aluBoi_shft_SRL_srl_16_U11 ( .B1(
        aluBoi_aluBoi_shft_SRL_srl_16_n1), .B2(
        aluBoi_aluBoi_shft_SRL_srl_16_n32), .C1(
        aluBoi_aluBoi_shft_SRL_srl_16_n4), .C2(
        aluBoi_aluBoi_shft_SRL_srl_16_n71), .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n180), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n124) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U10 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n108), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n3) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U9 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n6), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n5) );
  INV_X4 aluBoi_aluBoi_shft_SRL_srl_16_U8 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n9), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n8) );
  INV_X16 aluBoi_aluBoi_shft_SRL_srl_16_U7 ( .A(n6612), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n16) );
  INV_X16 aluBoi_aluBoi_shft_SRL_srl_16_U6 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n3), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n2) );
  INV_X8 aluBoi_aluBoi_shft_SRL_srl_16_U5 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n111), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n9) );
  INV_X16 aluBoi_aluBoi_shft_SRL_srl_16_U4 ( .A(
        aluBoi_aluBoi_shft_SRL_srl_16_n20), .ZN(
        aluBoi_aluBoi_shft_SRL_srl_16_n21) );
  INV_X2 aluBoi_aluBoi_shft_SRL_srl_16_U3 ( .A(aluBoi_aluBoi_shft_sraout[31]), 
        .ZN(aluBoi_aluBoi_shft_SRL_srl_16_n32) );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U65 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__1_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n6), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__1_) );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U64 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__0_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n16), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__0_) );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U63 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__1_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n16), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__1_) );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U62 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__2_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n16), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__2_) );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U61 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__3_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n16), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__3_) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U60 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__0_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n40) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U59 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__1_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n39) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U58 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__2_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n38) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U57 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__3_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n37) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U56 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__4_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n36) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U55 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__5_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n35) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U54 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__6_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n34) );
  NAND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U53 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__7_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n33) );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U52 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n40), .ZN(aluBoi_aluBoi_shft_sllout[0])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U51 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__10_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[10])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U50 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__11_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[11])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U49 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__12_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[12])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U48 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__13_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[13])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U47 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__14_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[14])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U46 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__15_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[15])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U45 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n39), .ZN(aluBoi_aluBoi_shft_sllout[1])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U44 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n38), .ZN(aluBoi_aluBoi_shft_sllout[2])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U43 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n37), .ZN(aluBoi_aluBoi_shft_sllout[3])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U42 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n36), .ZN(aluBoi_aluBoi_shft_sllout[4])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U41 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n35), .ZN(aluBoi_aluBoi_shft_sllout[5])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U40 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n34), .ZN(aluBoi_aluBoi_shft_sllout[6])
         );
  NOR2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U39 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_n23), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n33), .ZN(aluBoi_aluBoi_shft_sllout[7])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U38 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__8_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[8])
         );
  AND2_X1 aluBoi_aluBoi_shft_SLL_sll_7_U37 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__9_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_sllout[9])
         );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U36 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n39), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n32) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U35 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n38), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n31) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U34 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n40), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n30) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U33 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n37), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n29) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U32 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n35), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n28) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U31 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n34), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n27) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U30 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n36), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n26) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U29 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n33), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n25) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U28 ( .A(n6618), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n24) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U27 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n22) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U26 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n17), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n21) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U25 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n21), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n20) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U24 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n18), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n19) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U23 ( .A(n6616), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n18) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U22 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n18), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n17) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U21 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n16) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U20 ( .A(n6612), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n12) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U19 ( .A(n6612), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n11) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U18 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n1), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n8)
         );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U17 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n1), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n7)
         );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U16 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n1), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n6)
         );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U15 ( .A(n6606), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n2) );
  INV_X32 aluBoi_aluBoi_shft_SLL_sll_7_U14 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n2), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n1)
         );
  AND2_X4 aluBoi_aluBoi_shft_SLL_sll_7_U13 ( .A1(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__0_), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n6), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__0_) );
  AND2_X4 aluBoi_aluBoi_shft_SLL_sll_7_U12 ( .A1(net345751), .A2(
        aluBoi_aluBoi_shft_SLL_sll_7_n11), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__0_) );
  INV_X1 aluBoi_aluBoi_shft_SLL_sll_7_U11 ( .A(n6614), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n14) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U10 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n16), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n15) );
  INV_X4 aluBoi_aluBoi_shft_SLL_sll_7_U9 ( .A(aluBoi_aluBoi_shft_SLL_sll_7_n14), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n13) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U8 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n11), .ZN(
        aluBoi_aluBoi_shft_SLL_sll_7_n10) );
  INV_X8 aluBoi_aluBoi_shft_SLL_sll_7_U7 ( .A(aluBoi_aluBoi_shft_SLL_sll_7_n24), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n23) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U6 ( .A(aluBoi_aluBoi_shft_SLL_sll_7_n6), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n5) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U5 ( .A(aluBoi_aluBoi_shft_SLL_sll_7_n7), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n4) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U4 ( .A(aluBoi_aluBoi_shft_SLL_sll_7_n8), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n3) );
  INV_X16 aluBoi_aluBoi_shft_SLL_sll_7_U3 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_n12), .ZN(aluBoi_aluBoi_shft_SLL_sll_7_n9) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_1 ( .A(net368498), .B(net345751), 
        .S(n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__1_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_2 ( .A(net368502), .B(net368498), 
        .S(n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__2_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_3 ( .A(n13525), .B(net368502), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__3_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_4 ( .A(net377611), .B(n13525), .S(
        n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__4_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_5 ( .A(n6545), .B(net377611), .S(
        n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__5_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_6 ( .A(n6543), .B(n6545), .S(n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__6_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_7 ( .A(n6541), .B(n6543), .S(n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__7_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_8 ( .A(n5007), .B(n6541), .S(n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__8_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_9 ( .A(n13706), .B(n5007), .S(
        n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__9_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_10 ( .A(net368519), .B(n13706), 
        .S(n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__10_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_11 ( .A(n6539), .B(net368519), .S(
        n6612), .Z(aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__11_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_12 ( .A(n6537), .B(n6539), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__12_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_13 ( .A(n6535), .B(n6537), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__13_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_14 ( .A(n6533), .B(n6535), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__14_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_15 ( .A(n13527), .B(n6533), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__15_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_16 ( .A(n6529), .B(n13527), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__16_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_17 ( .A(n6527), .B(n6529), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__17_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_18 ( .A(n6525), .B(n6527), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__18_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_19 ( .A(n6523), .B(n6525), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__19_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_20 ( .A(n6521), .B(n6523), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__20_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_21 ( .A(n6519), .B(n6521), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__21_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_22 ( .A(net368572), .B(n6519), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n9), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__22_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_23 ( .A(net377607), .B(net368572), 
        .S(aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__23_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_24 ( .A(n5309), .B(net377607), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__24_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_25 ( .A(n6517), .B(n5309), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__25_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_26 ( .A(net368584), .B(n6517), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__26_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_27 ( .A(n6515), .B(net368584), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__27_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_28 ( .A(n6513), .B(n6515), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__28_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_29 ( .A(n6511), .B(n6513), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__29_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_30 ( .A(n6509), .B(n6511), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__30_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_0_31 ( .A(
        aluBoi_aluBoi_shft_sraout[31]), .B(n6509), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n10), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__31_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_2 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__2_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__0_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__2_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_3 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__3_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__1_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__3_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_4 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__4_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__2_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__4_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_5 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__5_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__3_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__5_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_6 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__6_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__4_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__6_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_7 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__7_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__5_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__7_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_8 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__8_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__6_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__8_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_9 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__9_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__7_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__9_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_10 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__10_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__8_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__10_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_11 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__11_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__9_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__11_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_12 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__12_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__10_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n3), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__12_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_13 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__13_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__11_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__13_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_14 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__14_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__12_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__14_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_15 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__15_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__13_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__15_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_16 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__16_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__14_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__16_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_17 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__17_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__15_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__17_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_18 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__18_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__16_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__18_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_19 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__19_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__17_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__19_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_20 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__20_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__18_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__20_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_21 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__21_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__19_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__21_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_22 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__22_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__20_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__22_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_23 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__23_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__21_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n4), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__23_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_24 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__24_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__22_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__24_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_25 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__25_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__23_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__25_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_26 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__26_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__24_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__26_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_27 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__27_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__25_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__27_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_28 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__28_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__26_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__28_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_29 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__29_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__27_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__29_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_30 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__30_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__28_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__30_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_1_31 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__31_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_1__29_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n5), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__31_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_4 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__4_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__0_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__4_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_5 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__5_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__1_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__5_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_6 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__6_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__2_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__6_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_7 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__7_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__3_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__7_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_8 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__8_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__4_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__8_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_9 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__9_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__5_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__9_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_10 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__10_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__6_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__10_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_11 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__11_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__7_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__11_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_12 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__12_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__8_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__12_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_13 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__13_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__9_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__13_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_14 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__14_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__10_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n13), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__14_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_15 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__15_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__11_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__15_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_16 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__16_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__12_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__16_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_17 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__17_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__13_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__17_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_18 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__18_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__14_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__18_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_19 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__19_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__15_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__19_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_20 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__20_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__16_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__20_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_21 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__21_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__17_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__21_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_22 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__22_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__18_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__22_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_23 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__23_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__19_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__23_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_24 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__24_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__20_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__24_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_25 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__25_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__21_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__25_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_26 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__26_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__22_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__26_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_27 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__27_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__23_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__27_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_28 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__28_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__24_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__28_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_29 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__29_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__25_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__29_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_30 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__30_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__26_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__30_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_2_31 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__31_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_2__27_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n15), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__31_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_8 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__8_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__0_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__8_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_9 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__9_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__1_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__9_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_10 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__10_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__2_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__10_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_11 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__11_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__3_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__11_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_12 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__12_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__4_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__12_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_13 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__13_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__5_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__13_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_14 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__14_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__6_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__14_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_15 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__15_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__7_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__15_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_16 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__16_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__8_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__16_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_17 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__17_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__9_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__17_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_18 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__18_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__10_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n19), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__18_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_19 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__19_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__11_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__19_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_20 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__20_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__12_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__20_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_21 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__21_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__13_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__21_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_22 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__22_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__14_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__22_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_23 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__23_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__15_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__23_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_24 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__24_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__16_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__24_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_25 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__25_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__17_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__25_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_26 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__26_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__18_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__26_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_27 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__27_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__19_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__27_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_28 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__28_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__20_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__28_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_29 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__29_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__21_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__29_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_30 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__30_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__22_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__30_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_3_31 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__31_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_3__23_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n20), .Z(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__31_) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_16 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__16_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n30), .S(aluBoi_aluBoi_shft_SLL_sll_7_n23), .Z(aluBoi_aluBoi_shft_sllout[16]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_17 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__17_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n32), .S(aluBoi_aluBoi_shft_SLL_sll_7_n23), .Z(aluBoi_aluBoi_shft_sllout[17]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_18 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__18_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n31), .S(aluBoi_aluBoi_shft_SLL_sll_7_n23), .Z(aluBoi_aluBoi_shft_sllout[18]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_19 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__19_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n29), .S(aluBoi_aluBoi_shft_SLL_sll_7_n23), .Z(aluBoi_aluBoi_shft_sllout[19]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_20 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__20_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n26), .S(aluBoi_aluBoi_shft_SLL_sll_7_n23), .Z(aluBoi_aluBoi_shft_sllout[20]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_21 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__21_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n28), .S(aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[21]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_22 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__22_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n27), .S(aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[22]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_23 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__23_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_n25), .S(aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[23]) );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_24 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__24_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__8_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[24])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_25 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__25_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__9_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[25])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_26 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__26_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__10_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[26])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_27 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__27_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__11_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[27])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_28 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__28_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__12_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[28])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_29 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__29_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__13_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[29])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_30 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__30_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__14_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[30])
         );
  MUX2_X2 aluBoi_aluBoi_shft_SLL_sll_7_M1_4_31 ( .A(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__31_), .B(
        aluBoi_aluBoi_shft_SLL_sll_7_ML_int_4__15_), .S(
        aluBoi_aluBoi_shft_SLL_sll_7_n22), .Z(aluBoi_aluBoi_shft_sllout[31])
         );
endmodule

